magic
tech scmos
timestamp 1385414349
<< pwell >>
rect -76 4 -48 14
rect -38 -15 132 -1
rect -38 -20 147 -15
rect -68 -39 147 -20
<< nwell >>
rect -76 22 132 42
rect -38 9 132 22
rect -79 -12 -48 -2
<< polysilicon >>
rect 48 56 52 60
rect -68 30 -64 32
rect -30 31 -26 52
rect -23 31 -19 44
rect -16 31 -12 33
rect 6 31 10 33
rect 34 31 38 44
rect 48 31 52 52
rect 82 31 86 44
rect 89 31 93 52
rect 121 48 125 60
rect 121 31 125 44
rect 135 31 139 52
rect -68 19 -64 26
rect -68 11 -64 15
rect -68 5 -64 7
rect -60 -5 -56 -3
rect -60 -13 -56 -9
rect -30 -16 -26 27
rect -23 -16 -19 27
rect -16 14 -12 27
rect -16 -16 -12 10
rect 6 14 10 27
rect 20 14 24 16
rect 6 -16 10 10
rect 20 6 24 10
rect 20 -2 24 2
rect 20 -8 24 -6
rect -60 -21 -56 -17
rect 34 -20 38 27
rect 48 -20 52 27
rect 82 -16 86 27
rect 89 -16 93 27
rect 107 20 111 22
rect 107 6 111 16
rect 107 -8 111 2
rect 107 -14 111 -12
rect 121 -16 125 27
rect 135 -16 139 27
rect -30 -22 -26 -20
rect -23 -22 -19 -20
rect -16 -22 -12 -20
rect 6 -22 10 -20
rect 82 -22 86 -20
rect 89 -22 93 -20
rect 121 -22 125 -20
rect 135 -22 139 -20
rect -60 -27 -56 -25
rect 34 -28 38 -24
rect 48 -28 52 -24
<< ndiffusion >>
rect -71 7 -68 11
rect -64 7 -61 11
rect 17 -6 20 -2
rect 24 -6 27 -2
rect -33 -20 -30 -16
rect -26 -20 -23 -16
rect -19 -20 -16 -16
rect -12 -20 -9 -16
rect 3 -20 6 -16
rect 10 -20 13 -16
rect 104 -12 107 -8
rect 111 -12 114 -8
rect 79 -20 82 -16
rect 86 -20 89 -16
rect 93 -20 96 -16
rect 118 -20 121 -16
rect 125 -20 128 -16
rect 132 -20 135 -16
rect 139 -20 142 -16
rect -63 -25 -60 -21
rect -56 -25 -53 -21
rect 30 -24 34 -20
rect 38 -24 41 -20
rect 45 -24 48 -20
rect 52 -24 55 -20
<< pdiffusion >>
rect -71 26 -68 30
rect -64 26 -61 30
rect -33 27 -30 31
rect -26 27 -23 31
rect -19 27 -16 31
rect -12 27 -9 31
rect 3 27 6 31
rect 10 27 14 31
rect 30 27 34 31
rect 38 27 41 31
rect 45 27 48 31
rect 52 27 55 31
rect 79 27 82 31
rect 86 27 89 31
rect 93 27 96 31
rect 118 27 121 31
rect 125 27 128 31
rect 132 27 135 31
rect 139 27 142 31
rect -63 -9 -60 -5
rect -56 -9 -53 -5
rect 17 10 20 14
rect 24 10 27 14
rect 104 16 107 20
rect 111 16 114 20
<< metal1 >>
rect -26 52 48 56
rect 52 52 89 56
rect 93 52 135 56
rect -19 44 34 48
rect 38 44 82 48
rect 86 44 121 48
rect -75 36 3 40
rect 20 36 146 40
rect -61 30 -57 36
rect -75 19 -71 26
rect -79 15 -71 19
rect -64 15 -61 19
rect -75 11 -71 15
rect -53 12 -49 36
rect -9 31 -5 36
rect -61 3 -57 7
rect -78 -1 -57 3
rect -1 31 3 36
rect 26 31 30 36
rect 55 31 59 36
rect 96 31 100 36
rect 114 31 118 36
rect 142 31 146 36
rect -37 6 -33 27
rect 14 23 18 27
rect 14 19 31 23
rect 27 14 31 19
rect 41 14 45 27
rect -12 10 -9 14
rect 3 10 6 14
rect 31 10 45 14
rect 13 6 17 10
rect 67 6 71 11
rect 75 6 79 27
rect 128 20 132 27
rect 118 16 132 20
rect 100 6 104 16
rect -78 -4 -74 -1
rect -53 -5 -49 6
rect -78 -33 -74 -10
rect -45 2 17 6
rect 24 2 104 6
rect 111 2 114 6
rect 118 2 150 6
rect -67 -21 -63 -9
rect -45 -13 -41 2
rect -56 -17 -41 -13
rect -37 -16 -33 2
rect 13 -2 17 2
rect 31 -6 45 -2
rect 27 -11 31 -6
rect 13 -15 31 -11
rect 13 -16 17 -15
rect -53 -33 -49 -25
rect -9 -33 -5 -20
rect 41 -20 45 -6
rect 75 -16 79 2
rect 100 -8 104 2
rect 118 -12 132 -8
rect 128 -16 132 -12
rect -1 -33 3 -20
rect 26 -33 30 -24
rect 55 -33 59 -24
rect 96 -33 100 -20
rect 114 -33 118 -20
rect 142 -33 146 -20
rect -78 -37 3 -33
rect 20 -37 146 -33
<< metal2 >>
rect -43 19 71 23
rect -57 15 -39 19
rect 67 15 71 19
rect -9 6 -5 10
rect -1 6 3 10
rect -9 2 63 6
rect 59 0 63 2
rect 114 0 118 2
rect 59 -4 118 0
rect -84 -17 -71 -13
rect -84 -39 -80 -17
rect -84 -43 49 -39
rect 45 -47 49 -43
<< ntransistor >>
rect -68 7 -64 11
rect 20 -6 24 -2
rect -30 -20 -26 -16
rect -23 -20 -19 -16
rect -16 -20 -12 -16
rect 6 -20 10 -16
rect 107 -12 111 -8
rect 82 -20 86 -16
rect 89 -20 93 -16
rect 121 -20 125 -16
rect 135 -20 139 -16
rect -60 -25 -56 -21
rect 34 -24 38 -20
rect 48 -24 52 -20
<< ptransistor >>
rect -68 26 -64 30
rect -30 27 -26 31
rect -23 27 -19 31
rect -16 27 -12 31
rect 6 27 10 31
rect 34 27 38 31
rect 48 27 52 31
rect 82 27 86 31
rect 89 27 93 31
rect 121 27 125 31
rect 135 27 139 31
rect -60 -9 -56 -5
rect 20 10 24 14
rect 107 16 111 20
<< polycontact >>
rect -30 52 -26 56
rect 48 52 52 56
rect -23 44 -19 48
rect 34 44 38 48
rect 89 52 93 56
rect 82 44 86 48
rect 121 44 125 48
rect 135 52 139 56
rect -68 15 -64 19
rect -60 -17 -56 -13
rect -16 10 -12 14
rect 6 10 10 14
rect 20 2 24 6
rect 107 2 111 6
<< ndcontact >>
rect -75 7 -71 11
rect -61 7 -57 11
rect 13 -6 17 -2
rect 27 -6 31 -2
rect -37 -20 -33 -16
rect -9 -20 -5 -16
rect -1 -20 3 -16
rect 13 -20 17 -16
rect 100 -12 104 -8
rect 114 -12 118 -8
rect 75 -20 79 -16
rect 96 -20 100 -16
rect 114 -20 118 -16
rect 128 -20 132 -16
rect 142 -20 146 -16
rect -67 -25 -63 -21
rect -53 -25 -49 -21
rect 26 -24 30 -20
rect 41 -24 45 -20
rect 55 -24 59 -20
<< pdcontact >>
rect -75 26 -71 30
rect -61 26 -57 30
rect -37 27 -33 31
rect -9 27 -5 31
rect -1 27 3 31
rect 14 27 18 31
rect 26 27 30 31
rect 41 27 45 31
rect 55 27 59 31
rect 75 27 79 31
rect 96 27 100 31
rect 114 27 118 31
rect 128 27 132 31
rect 142 27 146 31
rect -67 -9 -63 -5
rect -53 -9 -49 -5
rect 13 10 17 14
rect 27 10 31 14
rect 100 16 104 20
rect 114 16 118 20
<< m2contact >>
rect -61 15 -57 19
rect -9 10 -5 14
rect -1 10 3 14
rect 67 11 71 15
rect 114 2 118 6
rect -71 -17 -67 -13
<< psubstratepcontact >>
rect -53 6 -49 12
rect 3 -37 20 -33
<< nsubstratencontact >>
rect 3 36 20 40
rect -78 -10 -74 -4
<< labels >>
rlabel metal1 149 4 149 4 7 Cin
rlabel metal1 -78 17 -78 17 3 Cout
rlabel metal1 49 -36 49 -36 1 GND
rlabel metal2 47 -46 47 -46 1 S
rlabel metal1 49 39 49 39 5 Vdd
rlabel polysilicon 50 59 50 59 5 A
rlabel polysilicon 123 59 123 59 5 B
<< end >>
