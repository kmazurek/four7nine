magic
tech scmos
timestamp 1385331530
<< pwell >>
rect -17 -17 65 -7
rect -17 -47 40 -17
<< nwell >>
rect -17 3 25 21
<< polysilicon >>
rect -9 12 -5 24
rect 13 8 17 24
rect -9 -8 -5 8
rect -9 -24 -5 -12
rect 13 -16 17 4
rect 13 -32 17 -20
rect 36 -32 40 -4
rect 53 -8 57 -6
rect 53 -24 57 -12
rect 36 -38 40 -36
<< ndiffusion >>
rect -12 -12 -9 -8
rect -5 -12 -2 -8
rect 10 -20 13 -16
rect 17 -20 20 -16
rect 50 -12 53 -8
rect 57 -12 60 -8
rect 33 -36 36 -32
rect 40 -36 43 -32
<< pdiffusion >>
rect -12 8 -9 12
rect -5 8 -2 12
rect 10 4 13 8
rect 17 4 20 8
<< metal1 >>
rect -20 16 -1 20
rect 9 16 59 20
rect -16 12 -12 16
rect -2 0 2 8
rect 6 8 10 16
rect -2 -8 2 -4
rect 20 -8 24 4
rect 32 -4 36 0
rect 20 -12 46 -8
rect -16 -42 -12 -12
rect 20 -16 24 -12
rect -5 -28 -1 -24
rect 6 -42 10 -20
rect 60 -22 64 -12
rect 49 -28 53 -24
rect 60 -26 68 -22
rect 60 -32 64 -26
rect 17 -36 29 -32
rect 47 -36 64 -32
rect -20 -46 -12 -42
rect 6 -46 59 -42
<< metal2 >>
rect 2 -4 28 0
rect 3 -28 45 -24
<< ntransistor >>
rect -9 -12 -5 -8
rect 13 -20 17 -16
rect 53 -12 57 -8
rect 36 -36 40 -32
<< ptransistor >>
rect -9 8 -5 12
rect 13 4 17 8
<< polycontact >>
rect 36 -4 40 0
rect -9 -28 -5 -24
rect 53 -28 57 -24
rect 13 -36 17 -32
<< ndcontact >>
rect -16 -12 -12 -8
rect -2 -12 2 -8
rect 6 -20 10 -16
rect 20 -20 24 -16
rect 46 -12 50 -8
rect 60 -12 64 -8
rect 29 -36 33 -32
rect 43 -36 47 -32
<< pdcontact >>
rect -16 8 -12 12
rect -2 8 2 12
rect 6 4 10 8
rect 20 4 24 8
<< m2contact >>
rect -2 -4 2 0
rect 28 -4 32 0
rect -1 -28 3 -24
rect 45 -28 49 -24
<< psubstratepcontact >>
rect -12 -46 6 -42
<< nsubstratencontact >>
rect -1 16 9 20
<< labels >>
rlabel metal1 23 -45 23 -45 1 GND
rlabel metal1 23 19 23 19 5 Vdd
rlabel polysilicon -7 23 -7 23 5 In1
rlabel polysilicon 15 23 15 23 5 In2
rlabel metal1 67 -24 67 -24 7 Out
<< end >>
