magic
tech scmos
timestamp 1385900209
<< polysilicon >>
rect -43 26 -12 28
rect -43 19 -41 26
rect -20 19 -18 23
rect -8 19 -6 28
rect 1 21 16 23
rect 14 19 16 21
rect 25 19 27 22
rect 48 19 50 21
rect 100 19 102 26
rect 127 19 129 21
rect 138 19 140 21
rect 151 19 153 21
rect 178 19 180 22
rect -43 -7 -41 11
rect -43 -9 -38 -7
rect -34 -9 -32 -7
rect -20 -19 -18 11
rect -8 8 -6 11
rect 14 -10 16 11
rect 25 -10 27 11
rect 48 3 50 11
rect 35 1 50 3
rect 48 -11 50 1
rect 62 -4 64 5
rect 88 1 90 9
rect 88 -6 90 -3
rect 62 -11 64 -8
rect 48 -13 53 -11
rect 57 -13 59 -11
rect 100 -11 102 11
rect 127 1 129 11
rect 109 -1 129 1
rect 127 -10 129 -1
rect 138 -10 140 11
rect 151 1 153 11
rect 97 -13 105 -11
rect 109 -13 111 -11
rect 14 -17 16 -14
rect -51 -21 -15 -19
rect -11 -21 -9 -19
rect 25 -21 27 -14
rect 178 -11 180 11
rect 160 -13 183 -11
rect 187 -13 191 -11
rect 127 -17 129 -14
rect 138 -21 140 -14
<< ndiffusion >>
rect -38 -7 -34 -4
rect -38 -12 -34 -9
rect 11 -14 14 -10
rect 16 -14 18 -10
rect 22 -14 25 -10
rect 27 -14 31 -10
rect 85 -3 88 1
rect 90 -3 93 1
rect 57 -8 62 -4
rect 64 -8 67 -4
rect 53 -11 57 -8
rect 105 -11 109 -8
rect -15 -19 -11 -16
rect 53 -16 57 -13
rect 105 -16 109 -13
rect 124 -14 127 -10
rect 129 -14 131 -10
rect 135 -14 138 -10
rect 140 -14 144 -10
rect 183 -11 187 -8
rect 183 -16 187 -13
rect -15 -24 -11 -21
<< pdiffusion >>
rect -46 11 -43 19
rect -41 11 -38 19
rect -23 11 -20 19
rect -18 11 -15 19
rect -11 11 -8 19
rect -6 11 -3 19
rect 11 11 14 19
rect 16 11 25 19
rect 27 11 31 19
rect 45 11 48 19
rect 50 11 53 19
rect 97 11 100 19
rect 102 11 105 19
rect 124 11 127 19
rect 129 11 138 19
rect 140 11 144 19
rect 148 11 151 19
rect 153 11 156 19
rect 175 11 178 19
rect 180 11 183 19
<< metal1 >>
rect -55 55 192 63
rect -54 11 -50 55
rect -27 19 -23 55
rect -12 28 -8 34
rect -3 25 1 26
rect -3 19 1 21
rect 7 19 11 55
rect 41 19 45 55
rect -38 0 -34 11
rect -50 -9 -47 -5
rect -15 -12 -11 11
rect 31 -3 35 11
rect 18 -7 31 -3
rect 53 -4 57 11
rect 60 9 64 35
rect 18 -10 22 -7
rect 67 -4 71 26
rect 84 9 88 34
rect 93 19 97 55
rect 104 26 105 30
rect 120 19 124 55
rect 156 19 160 22
rect 80 -3 81 1
rect 93 -9 97 -3
rect 105 -4 109 11
rect 144 1 148 11
rect 163 5 167 34
rect 171 19 175 55
rect 157 1 167 5
rect 131 -3 148 1
rect 109 -8 111 -4
rect 131 -10 135 -3
rect 183 -4 187 11
rect 156 -9 160 -8
rect -38 -48 -34 -16
rect -15 -48 -11 -28
rect 7 -48 11 -14
rect 21 -25 25 -21
rect 31 -48 35 -14
rect 53 -48 57 -20
rect 105 -48 109 -20
rect 120 -48 124 -14
rect 134 -25 138 -21
rect 144 -48 148 -14
rect 183 -48 187 -20
rect -52 -56 192 -48
<< metal2 >>
rect -56 44 -38 48
rect -34 44 192 48
rect -56 34 -12 38
rect -8 35 60 38
rect 64 35 84 38
rect -8 34 84 35
rect 88 34 163 38
rect 167 34 192 38
rect -54 -5 -50 34
rect 1 26 67 30
rect 109 26 160 30
rect 35 -7 80 -3
rect 115 -8 156 -4
rect -50 -29 21 -25
rect 25 -29 134 -25
rect 138 -29 192 -25
<< ntransistor >>
rect -38 -9 -34 -7
rect 14 -14 16 -10
rect 25 -14 27 -10
rect 88 -3 90 1
rect 62 -8 64 -4
rect 53 -13 57 -11
rect 105 -13 109 -11
rect -15 -21 -11 -19
rect 127 -14 129 -10
rect 138 -14 140 -10
rect 183 -13 187 -11
<< ptransistor >>
rect -43 11 -41 19
rect -20 11 -18 19
rect -8 11 -6 19
rect 14 11 16 19
rect 25 11 27 19
rect 48 11 50 19
rect 100 11 102 19
rect 127 11 129 19
rect 138 11 140 19
rect 151 11 153 19
rect 178 11 180 19
<< polycontact >>
rect -12 24 -8 28
rect 100 26 104 30
rect -3 21 1 25
rect -47 -9 -43 -5
rect 35 3 39 7
rect 60 5 64 9
rect 84 5 88 9
rect 93 -13 97 -9
rect 109 1 113 5
rect 153 1 157 5
rect 21 -21 25 -17
rect 156 -13 160 -9
rect 134 -21 138 -17
<< ndcontact >>
rect -38 -4 -34 0
rect -38 -16 -34 -12
rect -15 -16 -11 -12
rect 7 -14 11 -10
rect 18 -14 22 -10
rect 31 -14 35 -10
rect 81 -3 85 1
rect 93 -3 97 1
rect 53 -8 57 -4
rect 67 -8 71 -4
rect 105 -8 109 -4
rect 53 -20 57 -16
rect 120 -14 124 -10
rect 131 -14 135 -10
rect 144 -14 148 -10
rect 183 -8 187 -4
rect 105 -20 109 -16
rect 183 -20 187 -16
rect -15 -28 -11 -24
<< pdcontact >>
rect -50 11 -46 19
rect -38 11 -34 19
rect -27 11 -23 19
rect -15 11 -11 19
rect -3 11 1 19
rect 7 11 11 19
rect 31 11 35 19
rect 41 11 45 19
rect 53 11 57 19
rect 93 11 97 19
rect 105 11 109 19
rect 120 11 124 19
rect 144 11 148 19
rect 156 11 160 19
rect 171 11 175 19
rect 183 11 187 19
<< m2contact >>
rect -38 44 -34 48
rect -12 34 -8 38
rect -3 26 1 30
rect 60 35 64 39
rect -54 -9 -50 -5
rect 31 -7 35 -3
rect 84 34 88 38
rect 67 26 71 30
rect 105 26 109 30
rect 163 34 167 38
rect 156 22 160 26
rect 76 -3 80 1
rect 111 -8 115 -4
rect 156 -8 160 -4
rect 21 -29 25 -25
rect 134 -29 138 -25
<< labels >>
rlabel metal1 183 0 187 4 3 Qout
rlabel metal1 -35 55 -32 63 7 Vdd
rlabel metal1 -34 -56 -30 -48 7 GND
rlabel metal2 -56 34 -52 38 7 clk
rlabel metal2 -56 44 -52 48 7 clkb
rlabel metal2 -50 -29 -46 -25 7 rst
rlabel polysilicon -51 -21 -47 -19 7 Din
<< end >>
