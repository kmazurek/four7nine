magic
tech scmos
timestamp 1385414154
<< polysilicon >>
rect -91 40 -89 55
rect -68 40 -66 60
rect -57 42 -43 44
rect -91 23 -89 36
rect -68 34 -66 36
rect -57 28 -55 42
rect -45 40 -43 42
rect -45 34 -43 36
rect -34 28 -32 60
rect -4 41 -2 56
rect 30 41 32 65
rect 50 41 52 56
rect 68 41 70 77
rect 78 41 80 43
rect 96 41 98 43
rect 107 42 138 44
rect -68 26 -55 28
rect -45 26 -32 28
rect -68 23 -66 26
rect -45 23 -43 26
rect -4 24 -2 37
rect 30 24 32 37
rect 50 35 52 37
rect 50 24 52 26
rect 68 24 70 37
rect 78 24 80 37
rect 96 24 98 37
rect -91 17 -89 19
rect -68 -4 -66 19
rect -45 15 -43 19
rect -4 18 -2 20
rect 30 18 32 20
rect 50 -4 52 20
rect 68 18 70 20
rect 78 18 80 20
rect 96 18 98 20
rect 107 -4 109 42
rect 116 41 118 42
rect 136 41 138 42
rect 116 34 118 37
rect 136 32 138 37
rect 116 24 118 27
rect 136 24 138 26
rect 116 19 118 20
rect 136 19 138 20
rect 144 19 146 60
rect 158 41 160 43
rect 183 41 185 43
rect 225 41 227 43
rect 248 41 250 60
rect 273 41 275 43
rect 283 41 285 73
rect 310 41 312 43
rect 158 24 160 37
rect 183 24 185 37
rect 225 24 227 37
rect 248 35 250 37
rect 248 24 250 27
rect 273 24 275 37
rect 283 24 285 37
rect 310 24 312 37
rect 116 17 146 19
rect 158 18 160 20
rect 183 18 185 20
rect 225 18 227 20
rect 248 -4 250 20
rect 273 18 275 20
rect 283 18 285 20
rect 310 18 312 20
<< ndiffusion >>
rect -92 19 -91 23
rect -89 19 -88 23
rect -69 19 -68 23
rect -66 19 -65 23
rect -46 19 -45 23
rect -43 19 -42 23
rect -5 20 -4 24
rect -2 20 -1 24
rect 29 20 30 24
rect 32 20 33 24
rect 49 20 50 24
rect 52 20 53 24
rect 67 20 68 24
rect 70 20 72 24
rect 76 20 78 24
rect 80 20 81 24
rect 95 20 96 24
rect 98 20 99 24
rect 115 20 116 24
rect 118 20 119 24
rect 135 20 136 24
rect 138 20 139 24
rect 157 20 158 24
rect 160 20 161 24
rect 182 20 183 24
rect 185 20 186 24
rect 224 20 225 24
rect 227 20 228 24
rect 247 20 248 24
rect 250 20 251 24
rect 272 20 273 24
rect 275 20 277 24
rect 281 20 283 24
rect 285 20 286 24
rect 309 20 310 24
rect 312 20 313 24
<< pdiffusion >>
rect -92 36 -91 40
rect -89 36 -88 40
rect -69 36 -68 40
rect -66 36 -65 40
rect -46 36 -45 40
rect -43 36 -42 40
rect -5 37 -4 41
rect -2 37 -1 41
rect 29 37 30 41
rect 32 37 33 41
rect 49 37 50 41
rect 52 37 53 41
rect 67 37 68 41
rect 70 37 78 41
rect 80 37 81 41
rect 95 37 96 41
rect 98 37 99 41
rect 115 37 116 41
rect 118 37 119 41
rect 135 37 136 41
rect 138 37 139 41
rect 157 37 158 41
rect 160 37 161 41
rect 182 37 183 41
rect 185 37 186 41
rect 224 37 225 41
rect 227 37 228 41
rect 247 37 248 41
rect 250 37 251 41
rect 272 37 273 41
rect 275 37 283 41
rect 285 37 286 41
rect 309 37 310 41
rect 312 37 313 41
<< metal1 >>
rect -9 73 70 77
rect 80 73 279 77
rect -9 65 26 69
rect 201 65 321 69
rect -76 56 -66 60
rect -60 56 -32 60
rect -26 56 -8 60
rect 2 56 49 60
rect 61 56 136 60
rect 144 56 250 60
rect 256 56 322 60
rect 29 45 75 49
rect 99 45 148 49
rect 203 45 261 49
rect 273 45 322 49
rect -1 44 322 45
rect -1 41 3 44
rect -96 23 -92 36
rect -73 23 -69 36
rect -65 23 -61 36
rect -50 23 -46 36
rect -42 23 -38 36
rect 25 41 29 44
rect 63 41 67 44
rect 91 41 95 44
rect 153 41 157 44
rect 178 41 182 44
rect 220 41 224 44
rect 268 41 272 44
rect 305 41 309 44
rect -9 24 -5 37
rect 33 31 37 37
rect 45 31 49 37
rect 33 27 49 31
rect 33 24 37 27
rect -1 8 3 20
rect 45 24 49 27
rect 53 34 57 37
rect 57 30 74 34
rect 81 31 85 37
rect 99 31 103 37
rect 111 31 115 37
rect 53 24 57 30
rect 85 27 92 31
rect 99 27 115 31
rect 99 24 103 27
rect 25 8 29 20
rect 63 8 67 20
rect 72 16 76 20
rect 81 8 85 20
rect 111 24 115 27
rect 119 31 123 37
rect 119 24 123 27
rect 131 31 135 37
rect 131 24 135 27
rect 139 31 143 37
rect 161 31 165 37
rect 186 31 190 37
rect 197 31 201 35
rect 228 31 232 37
rect 243 31 247 37
rect 139 27 147 31
rect 151 27 154 31
rect 161 27 169 31
rect 173 27 179 31
rect 186 27 201 31
rect 209 27 221 31
rect 228 27 247 31
rect 139 24 143 27
rect 161 24 165 27
rect 186 24 190 27
rect 228 24 232 27
rect 243 24 247 27
rect 251 31 255 37
rect 286 31 290 37
rect 251 27 269 31
rect 277 27 298 31
rect 302 27 306 31
rect 251 24 255 27
rect 277 24 281 27
rect 313 24 317 37
rect 91 8 95 20
rect 153 8 157 20
rect 178 8 182 20
rect 220 8 224 20
rect 268 8 272 20
rect 286 8 290 20
rect 305 8 309 20
rect 38 4 54 8
rect 101 4 148 8
rect 239 4 261 8
rect 290 4 299 8
rect -84 -4 -66 0
rect -60 -4 -13 0
rect -9 -4 40 0
rect 50 -4 109 0
rect 113 -4 244 0
rect 248 -4 322 0
<< metal2 >>
rect 53 51 123 55
rect 53 34 57 51
rect 119 31 123 51
rect 197 39 201 65
rect -13 0 -9 26
rect 81 16 85 27
rect 131 16 135 27
rect 173 27 205 31
rect 139 20 143 24
rect 76 12 135 16
rect 147 13 151 27
rect 298 13 302 27
rect 147 9 302 13
<< ntransistor >>
rect -91 19 -89 23
rect -68 19 -66 23
rect -45 19 -43 23
rect -4 20 -2 24
rect 30 20 32 24
rect 50 20 52 24
rect 68 20 70 24
rect 78 20 80 24
rect 96 20 98 24
rect 116 20 118 24
rect 136 20 138 24
rect 158 20 160 24
rect 183 20 185 24
rect 225 20 227 24
rect 248 20 250 24
rect 273 20 275 24
rect 283 20 285 24
rect 310 20 312 24
<< ptransistor >>
rect -91 36 -89 40
rect -68 36 -66 40
rect -45 36 -43 40
rect -4 37 -2 41
rect 30 37 32 41
rect 50 37 52 41
rect 68 37 70 41
rect 78 37 80 41
rect 96 37 98 41
rect 116 37 118 41
rect 136 37 138 41
rect 158 37 160 41
rect 183 37 185 41
rect 225 37 227 41
rect 248 37 250 41
rect 273 37 275 41
rect 283 37 285 41
rect 310 37 312 41
<< polycontact >>
rect 26 65 32 69
rect -66 56 -60 60
rect -32 56 -26 60
rect -8 56 2 60
rect 49 56 61 60
rect 70 73 80 77
rect 279 73 285 77
rect 136 56 144 60
rect 74 30 78 34
rect 92 27 96 31
rect -66 -4 -60 0
rect 40 -4 50 0
rect 250 56 256 60
rect 154 27 158 31
rect 179 27 183 31
rect 221 27 225 31
rect 269 27 273 31
rect 306 27 310 31
rect 109 -4 113 0
rect 244 -4 248 0
<< ndcontact >>
rect -96 19 -92 23
rect -88 19 -84 23
rect -73 19 -69 23
rect -65 19 -61 23
rect -50 19 -46 23
rect -42 19 -38 23
rect -9 20 -5 24
rect -1 20 3 24
rect 25 20 29 24
rect 33 20 37 24
rect 45 20 49 24
rect 53 20 57 24
rect 63 20 67 24
rect 72 20 76 24
rect 81 20 85 24
rect 91 20 95 24
rect 99 20 103 24
rect 111 20 115 24
rect 119 20 123 24
rect 131 20 135 24
rect 139 20 143 24
rect 153 20 157 24
rect 161 20 165 24
rect 178 20 182 24
rect 186 20 190 24
rect 220 20 224 24
rect 228 20 232 24
rect 243 20 247 24
rect 251 20 255 24
rect 268 20 272 24
rect 277 20 281 24
rect 286 20 290 24
rect 305 20 309 24
rect 313 20 317 24
<< pdcontact >>
rect -96 36 -92 40
rect -88 36 -84 40
rect -73 36 -69 40
rect -65 36 -61 40
rect -50 36 -46 40
rect -42 36 -38 40
rect -9 37 -5 41
rect -1 37 3 41
rect 25 37 29 41
rect 33 37 37 41
rect 45 37 49 41
rect 53 37 57 41
rect 63 37 67 41
rect 81 37 85 41
rect 91 37 95 41
rect 99 37 103 41
rect 111 37 115 41
rect 119 37 123 41
rect 131 37 135 41
rect 139 37 143 41
rect 153 37 157 41
rect 161 37 165 41
rect 178 37 182 41
rect 186 37 190 41
rect 220 37 224 41
rect 228 37 232 41
rect 243 37 247 41
rect 251 37 255 41
rect 268 37 272 41
rect 286 37 290 41
rect 305 37 309 41
rect 313 37 317 41
<< m2contact >>
rect 197 65 201 69
rect -13 26 -9 30
rect 53 30 57 34
rect 81 27 85 31
rect 72 12 76 16
rect 119 27 123 31
rect 131 27 135 31
rect 197 35 201 39
rect 147 27 151 31
rect 169 27 173 31
rect 205 27 209 31
rect 298 27 302 31
rect -13 -4 -9 0
<< psubstratepcontact >>
rect -1 4 38 8
rect 54 4 101 8
rect 148 4 239 8
rect 261 4 290 8
rect 299 4 328 8
<< nsubstratencontact >>
rect -1 45 29 49
rect 75 45 99 49
rect 148 45 203 49
rect 261 45 273 49
<< labels >>
rlabel metal1 41 46 42 47 1 Vdd
rlabel metal1 -7 66 -7 66 7 Din
rlabel metal1 -8 74 -8 74 7 rst
rlabel metal1 43 5 43 6 5 GND
rlabel metal1 106 29 106 29 1 no1
rlabel metal1 142 29 142 29 1 t2
rlabel metal1 40 29 40 29 1 n11
rlabel metal1 -6 -3 -6 -2 5 clkb
rlabel metal1 4 57 5 57 1 clk
rlabel m2contact 171 28 171 29 1 qbn
rlabel metal2 87 13 87 13 1 t2in
rlabel metal1 59 31 59 31 1 t1
rlabel metal1 316 28 316 28 3 Qoutb
rlabel metal1 319 67 320 67 3 Qout
<< end >>
