magic
tech scmos
timestamp 1386053849
use kris_bit_low_1bit  kris_bit_low_1bit_0
array 0 7 363 0 0 631
timestamp 1386053752
transform 1 0 -21 0 1 -4
box 21 4 384 635
<< end >>
