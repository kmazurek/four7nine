magic
tech scmos
timestamp 1385102351
<< pwell >>
rect -19 -28 112 5
<< nwell >>
rect -19 5 112 49
<< polysilicon >>
rect 0 35 2 37
rect 30 35 32 37
rect 51 35 53 37
rect 71 35 73 37
rect 91 35 93 37
rect 0 18 2 31
rect 11 18 13 20
rect 0 -9 2 14
rect 11 -1 13 14
rect 30 -1 32 31
rect 51 10 53 31
rect 71 28 73 31
rect 51 -1 53 6
rect 71 -1 73 24
rect 91 19 93 31
rect 91 -1 93 15
rect 11 -7 13 -5
rect 30 -11 32 -5
rect 51 -7 53 -5
rect 71 -7 73 -5
rect 91 -7 93 -5
rect 20 -13 32 -11
rect 0 -15 2 -13
<< ndiffusion >>
rect 9 -5 11 -1
rect 13 -5 15 -1
rect 27 -5 30 -1
rect 32 -5 35 -1
rect 48 -5 51 -1
rect 53 -5 56 -1
rect 68 -5 71 -1
rect 73 -5 76 -1
rect 88 -5 91 -1
rect 93 -5 96 -1
rect -2 -13 0 -9
rect 2 -13 4 -9
<< pdiffusion >>
rect -2 31 0 35
rect 2 31 4 35
rect 27 31 30 35
rect 32 31 35 35
rect 48 31 51 35
rect 53 31 56 35
rect 68 31 71 35
rect 73 31 76 35
rect 88 31 91 35
rect 93 31 96 35
<< metal1 >>
rect -19 41 19 48
rect 93 41 112 48
rect 23 35 27 41
rect 44 35 48 41
rect 64 35 68 41
rect 84 35 88 41
rect -9 31 -6 35
rect 8 31 19 35
rect 15 28 19 31
rect 15 24 22 28
rect -19 14 -2 18
rect 2 14 9 18
rect 13 14 15 18
rect 22 10 26 24
rect -19 6 9 10
rect -9 -3 -2 1
rect -6 -9 -2 -3
rect 5 -1 9 6
rect 15 6 26 10
rect 35 10 39 31
rect 56 10 60 31
rect 68 24 69 28
rect 35 6 49 10
rect 15 -1 19 6
rect 35 -1 39 6
rect 56 -1 60 6
rect 76 19 80 31
rect 96 28 100 31
rect 104 28 108 31
rect 96 24 108 28
rect 76 15 89 19
rect 76 -1 80 15
rect 96 -1 100 24
rect 107 14 112 18
rect 107 6 112 10
rect 8 -13 16 -9
rect 23 -20 27 -5
rect 44 -20 48 -5
rect 64 -20 68 -5
rect 84 -20 88 -5
rect -19 -27 18 -20
rect 92 -27 112 -20
<< metal2 >>
rect 104 35 108 49
rect -13 1 -9 31
rect 26 24 64 28
rect 19 14 103 18
rect 60 6 103 10
rect -13 -28 -9 -3
<< ntransistor >>
rect 11 -5 13 -1
rect 30 -5 32 -1
rect 51 -5 53 -1
rect 71 -5 73 -1
rect 91 -5 93 -1
rect 0 -13 2 -9
<< ptransistor >>
rect 0 31 2 35
rect 30 31 32 35
rect 51 31 53 35
rect 71 31 73 35
rect 91 31 93 35
<< polycontact >>
rect -2 14 2 18
rect 9 14 13 18
rect 69 24 73 28
rect 49 6 53 10
rect 89 15 93 19
rect 16 -13 20 -9
<< ndcontact >>
rect 5 -5 9 -1
rect 15 -5 19 -1
rect 23 -5 27 -1
rect 35 -5 39 -1
rect 44 -5 48 -1
rect 56 -5 60 -1
rect 64 -5 68 -1
rect 76 -5 80 -1
rect 84 -5 88 -1
rect 96 -5 100 -1
rect -6 -13 -2 -9
rect 4 -13 8 -9
<< pdcontact >>
rect -6 31 -2 35
rect 4 31 8 35
rect 23 31 27 35
rect 35 31 39 35
rect 44 31 48 35
rect 56 31 60 35
rect 64 31 68 35
rect 76 31 80 35
rect 84 31 88 35
rect 96 31 100 35
<< m2contact >>
rect -13 31 -9 35
rect 22 24 26 28
rect 15 14 19 18
rect -13 -3 -9 1
rect 64 24 68 28
rect 56 6 60 10
rect 104 31 108 35
rect 103 14 107 18
rect 103 6 107 10
<< psubstratepcontact >>
rect 18 -27 92 -20
<< nsubstratencontact >>
rect 19 41 93 48
<< labels >>
rlabel metal1 -19 6 -7 10 7 inbit
rlabel metal1 -19 14 -7 18 7 shift
rlabel metal1 105 6 112 10 3 inbit_next
rlabel metal1 103 14 112 18 3 shift
rlabel metal2 -13 -28 -9 -28 5 shiftbit_in
rlabel metal2 104 49 108 49 1 shiftbit_out
rlabel metal1 -10 44 -10 44 5 Vdd
rlabel metal1 -7 -24 -7 -24 1 GND
<< end >>
