magic
tech scmos
timestamp 1385602182
<< pwell >>
rect -51 91 240 127
<< nwell >>
rect -51 127 240 173
<< polysilicon >>
rect -41 137 -39 139
rect -31 137 -29 151
rect -13 137 -11 140
rect 11 137 13 152
rect 28 137 30 161
rect 44 137 46 152
rect 62 137 64 139
rect 72 137 74 168
rect 130 140 132 156
rect 90 137 92 139
rect 110 138 132 140
rect 110 137 112 138
rect 130 137 132 138
rect 152 137 154 139
rect 177 137 179 139
rect 201 137 203 139
rect 211 137 213 168
rect 227 137 229 156
rect -41 120 -39 133
rect -31 120 -29 133
rect -13 120 -11 133
rect 11 120 13 133
rect 28 120 30 133
rect 44 131 46 133
rect 44 120 46 122
rect 62 120 64 133
rect 72 120 74 133
rect 90 120 92 133
rect 110 130 112 133
rect 130 128 132 133
rect 110 120 112 123
rect 130 120 132 122
rect 152 120 154 133
rect 177 120 179 133
rect 201 120 203 133
rect 211 120 213 133
rect 227 131 229 133
rect 227 120 229 123
rect -41 114 -39 116
rect -31 114 -29 116
rect -13 114 -11 116
rect 11 114 13 116
rect 28 114 30 116
rect 44 92 46 116
rect 62 114 64 116
rect 72 114 74 116
rect 90 114 92 116
rect 110 115 112 116
rect 130 115 132 116
rect 110 113 132 115
rect 152 114 154 116
rect 177 114 179 116
rect 110 92 112 113
rect 201 111 203 116
rect 211 114 213 116
rect 193 107 203 111
rect 227 92 229 116
<< ndiffusion >>
rect -42 116 -41 120
rect -39 116 -31 120
rect -29 116 -28 120
rect -14 116 -13 120
rect -11 116 -10 120
rect 10 116 11 120
rect 13 116 14 120
rect 27 116 28 120
rect 30 116 31 120
rect 43 116 44 120
rect 46 116 47 120
rect 61 116 62 120
rect 64 116 66 120
rect 70 116 72 120
rect 74 116 75 120
rect 89 116 90 120
rect 92 116 93 120
rect 109 116 110 120
rect 112 116 113 120
rect 129 116 130 120
rect 132 116 133 120
rect 151 116 152 120
rect 154 116 155 120
rect 176 116 177 120
rect 179 116 180 120
rect 200 116 201 120
rect 203 116 205 120
rect 209 116 211 120
rect 213 116 214 120
rect 226 116 227 120
rect 229 116 230 120
<< pdiffusion >>
rect -42 133 -41 137
rect -39 133 -37 137
rect -33 133 -31 137
rect -29 133 -28 137
rect -14 133 -13 137
rect -11 133 -10 137
rect 10 133 11 137
rect 13 133 14 137
rect 27 133 28 137
rect 30 133 31 137
rect 43 133 44 137
rect 46 133 47 137
rect 61 133 62 137
rect 64 133 72 137
rect 74 133 75 137
rect 89 133 90 137
rect 92 133 93 137
rect 109 133 110 137
rect 112 133 113 137
rect 129 133 130 137
rect 132 133 133 137
rect 151 133 152 137
rect 154 133 155 137
rect 176 133 177 137
rect 179 133 180 137
rect 200 133 201 137
rect 203 133 211 137
rect 213 133 214 137
rect 226 133 227 137
rect 229 133 230 137
<< metal1 >>
rect -51 168 64 172
rect 74 168 207 172
rect 213 168 240 172
rect -51 161 24 165
rect -2 152 11 156
rect 17 152 43 156
rect 55 152 132 156
rect 140 152 229 156
rect -51 141 -28 145
rect 2 141 14 145
rect 27 141 142 145
rect 201 141 240 145
rect -46 140 240 141
rect -46 137 -42 140
rect -28 137 -24 140
rect -18 137 -14 140
rect 14 137 18 140
rect -37 129 -33 133
rect -51 125 -45 129
rect -37 125 -17 129
rect -28 120 -24 125
rect -10 120 -6 133
rect 23 137 27 140
rect 57 137 61 140
rect 85 137 89 140
rect 147 137 151 140
rect 172 137 176 140
rect 196 137 200 140
rect 6 120 10 133
rect 31 127 35 133
rect 39 127 43 133
rect 31 123 43 127
rect 31 120 35 123
rect -46 104 -42 116
rect -18 104 -14 116
rect 14 104 18 116
rect 39 120 43 123
rect 47 130 51 133
rect 51 126 58 130
rect 75 127 79 133
rect 93 127 97 133
rect 105 127 109 133
rect 47 120 51 126
rect 66 123 80 127
rect 84 123 86 127
rect 93 123 109 127
rect 66 120 70 123
rect 93 120 97 123
rect 23 104 27 116
rect 57 104 61 116
rect 75 104 79 116
rect 105 120 109 123
rect 113 127 117 133
rect 113 120 117 123
rect 125 127 129 133
rect 125 120 129 123
rect 133 127 137 133
rect 155 127 159 133
rect 180 127 184 133
rect 187 127 191 131
rect 214 127 218 133
rect 222 127 226 133
rect 133 123 141 127
rect 145 123 148 127
rect 155 123 173 127
rect 180 123 191 127
rect 205 123 226 127
rect 230 127 234 133
rect 133 120 137 123
rect 155 120 159 123
rect 85 104 89 116
rect 147 104 151 116
rect 163 111 167 123
rect 180 120 184 123
rect 205 120 209 123
rect 222 120 226 123
rect 172 104 176 116
rect 184 107 189 111
rect 196 104 200 116
rect 214 104 218 116
rect -51 100 -47 104
rect -8 100 14 104
rect 36 100 48 104
rect 95 100 163 104
rect 203 100 240 104
rect 6 92 36 96
rect 44 92 106 96
rect 110 92 223 96
<< metal2 >>
rect 187 159 240 163
rect -6 128 -2 152
rect 47 147 117 151
rect 47 130 51 147
rect 113 127 117 147
rect 187 135 191 159
rect 2 96 6 122
rect 80 112 84 123
rect 121 112 125 127
rect 133 116 137 120
rect 80 108 125 112
rect 141 100 145 123
rect 167 107 180 111
rect 230 100 234 123
rect 141 96 234 100
<< ntransistor >>
rect -41 116 -39 120
rect -31 116 -29 120
rect -13 116 -11 120
rect 11 116 13 120
rect 28 116 30 120
rect 44 116 46 120
rect 62 116 64 120
rect 72 116 74 120
rect 90 116 92 120
rect 110 116 112 120
rect 130 116 132 120
rect 152 116 154 120
rect 177 116 179 120
rect 201 116 203 120
rect 211 116 213 120
rect 227 116 229 120
<< ptransistor >>
rect -41 133 -39 137
rect -31 133 -29 137
rect -13 133 -11 137
rect 11 133 13 137
rect 28 133 30 137
rect 44 133 46 137
rect 62 133 64 137
rect 72 133 74 137
rect 90 133 92 137
rect 110 133 112 137
rect 130 133 132 137
rect 152 133 154 137
rect 177 133 179 137
rect 201 133 203 137
rect 211 133 213 137
rect 227 133 229 137
<< polycontact >>
rect 64 168 74 172
rect 207 168 213 172
rect 24 161 30 165
rect 11 152 17 156
rect 43 152 55 156
rect 132 152 140 156
rect 229 152 235 156
rect -45 125 -41 129
rect -17 125 -13 129
rect 58 126 62 130
rect 86 123 90 127
rect 148 123 152 127
rect 173 123 177 127
rect 36 92 44 96
rect 106 92 110 96
rect 189 107 193 111
rect 223 92 227 96
<< ndcontact >>
rect -46 116 -42 120
rect -28 116 -24 120
rect -18 116 -14 120
rect -10 116 -6 120
rect 6 116 10 120
rect 14 116 18 120
rect 23 116 27 120
rect 31 116 35 120
rect 39 116 43 120
rect 47 116 51 120
rect 57 116 61 120
rect 66 116 70 120
rect 75 116 79 120
rect 85 116 89 120
rect 93 116 97 120
rect 105 116 109 120
rect 113 116 117 120
rect 125 116 129 120
rect 133 116 137 120
rect 147 116 151 120
rect 155 116 159 120
rect 172 116 176 120
rect 180 116 184 120
rect 196 116 200 120
rect 205 116 209 120
rect 214 116 218 120
rect 222 116 226 120
rect 230 116 234 120
<< pdcontact >>
rect -46 133 -42 137
rect -37 133 -33 137
rect -28 133 -24 137
rect -18 133 -14 137
rect -10 133 -6 137
rect 6 133 10 137
rect 14 133 18 137
rect 23 133 27 137
rect 31 133 35 137
rect 39 133 43 137
rect 47 133 51 137
rect 57 133 61 137
rect 75 133 79 137
rect 85 133 89 137
rect 93 133 97 137
rect 105 133 109 137
rect 113 133 117 137
rect 125 133 129 137
rect 133 133 137 137
rect 147 133 151 137
rect 155 133 159 137
rect 172 133 176 137
rect 180 133 184 137
rect 196 133 200 137
rect 214 133 218 137
rect 222 133 226 137
rect 230 133 234 137
<< m2contact >>
rect -6 152 -2 156
rect -6 124 -2 128
rect 2 122 6 126
rect 47 126 51 130
rect 80 123 84 127
rect 113 123 117 127
rect 125 123 129 127
rect 187 131 191 135
rect 141 123 145 127
rect 230 123 234 127
rect 163 107 167 111
rect 180 107 184 111
rect 2 92 6 96
<< psubstratepcontact >>
rect -47 100 -8 104
rect 14 100 36 104
rect 48 100 95 104
rect 163 100 203 104
<< nsubstratencontact >>
rect -28 141 2 145
rect 14 141 27 145
rect 142 141 201 145
<< labels >>
rlabel metal1 -2 163 -2 163 7 D
rlabel metal1 220 155 220 155 5 clk
rlabel metal1 36 144 36 144 5 Vdd
rlabel metal1 39 101 39 101 1 GND
rlabel metal1 -51 125 -51 129 7 load
rlabel metal1 2 153 2 154 1 clk1
rlabel polysilicon -30 150 -30 150 1 clk
rlabel metal2 239 161 239 161 3 Q
rlabel metal1 -51 161 -51 165 7 D
rlabel metal1 10 93 11 93 1 clkb
rlabel metal1 -51 100 -51 104 3 GND
rlabel metal1 240 100 240 104 7 GND
rlabel metal1 -51 168 -51 172 7 rst
rlabel metal1 239 170 239 170 3 rst
rlabel metal1 240 140 240 145 7 Vdd
<< end >>
