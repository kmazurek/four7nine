magic
tech scmos
timestamp 1386032703
<< pwell >>
rect 227 -656 266 -649
rect 220 -662 266 -656
rect 187 -680 271 -662
<< polysilicon >>
rect 7 39 9 142
rect 7 37 38 39
<< metal1 >>
rect -41 113 321 121
rect 262 58 272 62
rect 262 22 266 58
rect -41 2 322 10
rect -41 -7 -27 -3
rect -41 -15 -27 -11
rect -41 -35 -27 -31
rect 31 -35 101 -31
rect -41 -77 -27 -73
rect 35 -77 39 -73
rect 43 -77 48 -73
rect -41 -85 -27 -81
rect 35 -85 48 -81
rect -41 -93 -27 -89
rect 35 -93 48 -89
rect -41 -101 -27 -97
rect 35 -101 48 -97
rect -41 -109 -27 -105
rect 35 -109 48 -105
rect -41 -117 -27 -113
rect 35 -117 48 -113
rect -41 -125 -27 -121
rect 35 -125 48 -121
rect -41 -133 -27 -129
rect 35 -133 48 -129
rect -41 -141 -27 -137
rect 35 -141 48 -137
rect -41 -165 -27 -161
rect 19 -195 23 -186
rect -41 -199 23 -195
rect 53 -256 159 -252
rect -41 -265 -27 -261
rect -41 -273 -27 -269
rect -41 -281 -27 -277
rect -41 -288 -27 -284
rect -41 -296 -27 -292
rect -41 -304 -27 -300
rect -41 -312 -27 -308
rect -41 -320 -27 -316
rect -41 -328 -27 -324
rect -41 -336 -27 -332
rect -41 -344 -27 -340
rect -41 -352 -27 -348
rect -41 -360 -27 -356
rect -41 -368 -27 -364
rect -41 -376 -27 -372
rect -41 -384 -27 -380
rect -41 -392 -27 -388
rect -41 -400 -27 -396
rect -41 -408 -27 -404
rect -41 -415 -27 -411
rect -41 -423 -27 -419
rect -41 -431 -27 -427
rect -41 -439 -27 -435
rect -41 -447 -27 -443
rect -41 -455 -27 -451
rect -41 -463 -27 -459
rect -41 -471 -27 -467
rect -41 -479 -27 -475
rect -41 -487 -27 -483
rect -41 -495 -27 -491
rect -41 -503 -27 -499
rect -41 -511 -27 -507
rect -41 -522 -38 -518
rect -41 -531 -34 -527
rect -41 -539 -38 -535
rect -35 -664 -28 -661
rect -35 -668 62 -664
rect 69 -668 75 -664
rect 88 -733 322 -729
rect 86 -763 216 -756
rect 223 -763 322 -756
<< metal2 >>
rect -41 92 46 96
rect 271 92 322 96
rect -41 29 46 33
rect 271 29 322 33
rect 39 -198 43 -77
rect 177 -161 181 -15
rect 241 -234 245 -3
rect 262 -11 266 18
rect 159 -252 163 -251
rect -33 -646 -29 -635
rect -33 -650 85 -646
rect 62 -688 69 -668
rect 81 -692 85 -650
rect 216 -756 223 -617
<< polycontact >>
rect 101 -35 105 -31
rect 162 -85 166 -81
rect 49 -256 53 -252
rect 31 -265 35 -261
rect 67 -273 71 -269
<< m2contact >>
rect 262 18 266 22
rect 177 -15 181 -11
rect 262 -15 266 -11
rect 39 -77 43 -73
rect 177 -165 181 -161
rect 39 -202 43 -198
rect 241 -238 245 -234
rect 159 -256 163 -252
rect 216 -617 223 -613
rect -33 -635 -29 -631
rect 62 -668 69 -661
rect 62 -695 69 -688
rect 216 -763 223 -756
use reg2_na  reg2_na_0
timestamp 1385921827
transform 1 0 89 0 1 58
box -59 -56 193 63
use add1_flat_first  add1_flat_first_0
timestamp 1385746031
transform 1 0 -248 0 1 -318
box 278 66 516 315
use mux1  mux1_0
timestamp 1385747650
transform 1 0 87 0 1 -681
box -128 -18 235 678
use shift1  shift1_0
timestamp 1385746524
transform -1 0 71 0 -1 -715
box -19 -28 112 49
<< labels >>
rlabel metal1 37 -34 37 -34 1 Qout
rlabel metal2 -32 -647 -31 -647 3 shiftbit_in
<< end >>
