magic
tech scmos
timestamp 1385668156
<< pwell >>
rect 227 -656 266 -649
rect 220 -662 266 -656
rect 187 -680 271 -662
<< metal1 >>
rect 295 77 361 81
rect 295 69 361 73
rect 89 26 93 34
rect 354 33 362 37
rect 93 -35 195 -31
rect -32 -77 124 -73
rect 129 -77 142 -73
rect -32 -85 124 -81
rect 129 -85 142 -81
rect -32 -93 124 -89
rect 129 -93 142 -89
rect -32 -101 124 -97
rect 129 -101 142 -97
rect -32 -109 124 -105
rect 129 -109 142 -105
rect -32 -117 124 -113
rect 129 -117 142 -113
rect -32 -125 124 -121
rect 129 -125 142 -121
rect -32 -133 124 -129
rect 129 -133 142 -129
rect -32 -141 124 -137
rect 129 -141 142 -137
rect 53 -256 257 -252
rect -31 -668 62 -664
rect 69 -668 75 -664
<< metal2 >>
rect 89 -31 93 22
rect 311 4 315 8
rect 311 0 339 4
rect 335 -234 339 0
rect 356 -11 360 49
rect -40 -646 -36 -635
rect -40 -650 85 -646
rect 62 -688 69 -668
rect 81 -692 85 -650
<< polycontact >>
rect 350 33 354 37
rect 195 -35 199 -31
rect 49 -256 53 -252
<< m2contact >>
rect 356 49 360 53
rect 89 22 93 26
rect 311 8 315 12
rect 356 -15 360 -11
rect 89 -35 93 -31
rect 335 -238 339 -234
rect 253 -252 257 -248
rect -40 -635 -36 -631
rect 62 -668 69 -661
rect 62 -695 69 -688
use add1_flat_first  add1_flat_first_0
timestamp 1385598647
transform 1 0 -154 0 1 -318
box 278 66 516 315
use mux1  mux1_0
timestamp 1385599424
transform 1 0 87 0 1 -681
box -127 -6 275 678
use shift1  shift1_0
timestamp 1385102351
transform -1 0 72 0 -1 -715
box -19 -28 112 49
<< labels >>
rlabel metal1 362 33 362 37 3 load
rlabel space -37 9 365 88 1 REGISTER_GOES_HERE
rlabel metal2 -39 -647 -38 -647 3 shiftbit_in
rlabel space -51 -884 326 -768 1 REGISTER_GOES_HERE
<< end >>
