magic
tech scmos
timestamp 1385597418
<< pwell >>
rect -150 -113 -94 -99
rect -149 -125 -94 -113
rect -150 -197 -94 -175
rect -58 -197 -24 -179
<< nwell >>
rect -150 -89 -94 -57
rect -150 -165 -94 -143
rect -58 -157 -35 -143
<< polysilicon >>
rect -120 -76 -116 -74
rect -106 -76 -102 -74
rect -142 -84 -138 -82
rect -142 -92 -138 -88
rect -142 -100 -138 -96
rect -120 -100 -116 -80
rect -142 -106 -138 -104
rect -120 -108 -116 -104
rect -106 -87 -102 -80
rect -106 -108 -102 -91
rect -94 -104 -83 -100
rect -120 -114 -116 -112
rect -106 -114 -102 -112
rect -95 -124 -63 -120
rect -120 -152 -116 -150
rect -106 -152 -102 -150
rect -50 -152 -46 -150
rect -142 -160 -138 -158
rect -142 -168 -138 -164
rect -142 -176 -138 -172
rect -120 -176 -116 -156
rect -142 -182 -138 -180
rect -120 -184 -116 -180
rect -106 -163 -102 -156
rect -106 -184 -102 -167
rect -50 -168 -46 -156
rect -50 -184 -46 -172
rect -120 -190 -116 -188
rect -106 -190 -102 -188
rect -50 -190 -46 -188
<< ndiffusion >>
rect -145 -104 -142 -100
rect -138 -104 -135 -100
rect -123 -112 -120 -108
rect -116 -112 -106 -108
rect -102 -112 -99 -108
rect -145 -180 -142 -176
rect -138 -180 -135 -176
rect -123 -188 -120 -184
rect -116 -188 -106 -184
rect -102 -188 -99 -184
rect -53 -188 -50 -184
rect -46 -188 -43 -184
<< pdiffusion >>
rect -123 -80 -120 -76
rect -116 -80 -113 -76
rect -109 -80 -106 -76
rect -102 -80 -99 -76
rect -145 -88 -142 -84
rect -138 -88 -135 -84
rect -123 -156 -120 -152
rect -116 -156 -113 -152
rect -109 -156 -106 -152
rect -102 -156 -99 -152
rect -53 -156 -50 -152
rect -46 -156 -43 -152
rect -145 -164 -142 -160
rect -138 -164 -135 -160
<< metal1 >>
rect -21 -45 78 -41
rect -21 -50 -17 -45
rect 5 -54 33 -50
rect -150 -62 -149 -58
rect -136 -62 -90 -58
rect -86 -62 -63 -58
rect -135 -84 -131 -62
rect -127 -76 -123 -62
rect -99 -76 -95 -62
rect 33 -78 37 -54
rect -149 -92 -145 -88
rect -113 -92 -109 -80
rect -102 -91 -86 -87
rect -157 -96 -145 -92
rect -138 -96 -109 -92
rect -149 -100 -145 -96
rect -135 -120 -131 -104
rect -127 -108 -123 -96
rect -116 -104 -98 -100
rect -99 -120 -95 -112
rect -150 -124 -149 -120
rect -136 -124 -99 -120
rect -90 -128 -86 -91
rect -79 -104 -75 -100
rect 33 -128 37 -82
rect -90 -132 33 -128
rect 55 -102 59 -45
rect 66 -54 78 -50
rect 55 -106 78 -102
rect 55 -128 59 -106
rect 59 -132 78 -128
rect -157 -140 -57 -136
rect -35 -140 -9 -136
rect -35 -144 -31 -140
rect -150 -148 -149 -144
rect -136 -148 -90 -144
rect -86 -148 -47 -144
rect -36 -148 -31 -144
rect -135 -160 -131 -148
rect -127 -152 -123 -148
rect -99 -152 -95 -148
rect -43 -152 -39 -148
rect -149 -168 -145 -164
rect -113 -168 -109 -156
rect -102 -167 -75 -163
rect -157 -172 -145 -168
rect -138 -172 -109 -168
rect -57 -168 -53 -156
rect -46 -172 -18 -168
rect -149 -176 -145 -172
rect -135 -192 -131 -180
rect -127 -184 -123 -172
rect -116 -180 -112 -176
rect -99 -192 -95 -188
rect -150 -196 -149 -192
rect -136 -196 -94 -192
rect -81 -206 -77 -180
rect -57 -184 -53 -172
rect -22 -182 -18 -172
rect -43 -192 -39 -188
rect -69 -196 -65 -192
rect -61 -196 -57 -192
rect -46 -196 -20 -192
rect -24 -198 -20 -196
rect -24 -202 -9 -198
rect 74 -206 78 -132
rect -81 -210 78 -206
<< metal2 >>
rect 37 -54 62 -50
rect -90 -144 -86 -62
rect 37 -82 78 -78
rect -75 -163 -71 -104
rect -55 -128 -51 -124
rect -65 -132 -51 -128
rect -108 -180 -81 -176
rect -65 -192 -61 -132
rect -57 -168 -53 -140
rect -90 -196 -73 -192
<< ntransistor >>
rect -142 -104 -138 -100
rect -120 -112 -116 -108
rect -106 -112 -102 -108
rect -142 -180 -138 -176
rect -120 -188 -116 -184
rect -106 -188 -102 -184
rect -50 -188 -46 -184
<< ptransistor >>
rect -120 -80 -116 -76
rect -106 -80 -102 -76
rect -142 -88 -138 -84
rect -120 -156 -116 -152
rect -106 -156 -102 -152
rect -50 -156 -46 -152
rect -142 -164 -138 -160
<< polycontact >>
rect -21 -54 -17 -50
rect 1 -54 5 -50
rect -142 -96 -138 -92
rect -120 -104 -116 -100
rect -106 -91 -102 -87
rect -98 -104 -94 -100
rect -83 -104 -79 -100
rect -99 -124 -95 -120
rect -63 -124 -59 -120
rect 33 -132 37 -128
rect 55 -132 59 -128
rect -142 -172 -138 -168
rect -120 -180 -116 -176
rect -106 -167 -102 -163
rect -50 -172 -46 -168
<< ndcontact >>
rect -149 -104 -145 -100
rect -135 -104 -131 -100
rect -127 -112 -123 -108
rect -99 -112 -95 -108
rect -149 -180 -145 -176
rect -135 -180 -131 -176
rect -127 -188 -123 -184
rect -99 -188 -95 -184
rect -57 -188 -53 -184
rect -43 -188 -39 -184
<< pdcontact >>
rect -127 -80 -123 -76
rect -113 -80 -109 -76
rect -99 -80 -95 -76
rect -149 -88 -145 -84
rect -135 -88 -131 -84
rect -127 -156 -123 -152
rect -113 -156 -109 -152
rect -99 -156 -95 -152
rect -57 -156 -53 -152
rect -43 -156 -39 -152
rect -149 -164 -145 -160
rect -135 -164 -131 -160
<< m2contact >>
rect 33 -54 37 -50
rect -90 -62 -86 -58
rect 33 -82 37 -78
rect -75 -104 -71 -100
rect -55 -124 -51 -120
rect 62 -54 66 -50
rect -57 -140 -53 -136
rect -90 -148 -86 -144
rect -75 -167 -71 -163
rect -57 -172 -53 -168
rect -112 -180 -108 -176
rect -81 -180 -77 -176
rect -94 -196 -90 -192
rect -73 -196 -69 -192
rect -65 -196 -61 -192
<< psubstratepcontact >>
rect -149 -124 -136 -120
rect -149 -196 -136 -192
rect -57 -196 -46 -192
<< nsubstratencontact >>
rect -149 -62 -136 -58
rect -149 -148 -136 -144
rect -47 -148 -36 -144
use XOR  XOR_0
timestamp 1385331530
transform -1 0 -4 0 1 -78
box -20 -47 68 24
use XOR  XOR_1
timestamp 1385331530
transform -1 0 50 0 1 -156
box -20 -47 68 24
<< labels >>
rlabel metal1 -156 -138 -156 -138 3 Out00
rlabel metal1 -82 -59 -82 -59 5 Vdd
rlabel metal1 -83 -145 -83 -145 5 Vdd
rlabel metal1 -156 -94 -156 -94 3 Out10
rlabel metal1 -156 -170 -156 -170 3 Out01
rlabel metal1 -65 -195 -65 -195 1 GND
rlabel metal2 77 -80 77 -80 7 Sel0
rlabel metal1 77 -104 77 -104 7 Sel1
rlabel metal1 78 -54 78 -50 7 sel0
rlabel metal1 78 -45 78 -41 6 sel1
<< end >>
