magic
tech scmos
timestamp 1386053941
use data_high_final  data_high_final_0
timestamp 1386053173
transform 1 0 -653 0 1 279
box 653 -279 3557 753
use data_low_final  data_low_final_0
timestamp 1386053849
transform 1 0 2904 0 1 0
box 0 0 2904 631
<< end >>
