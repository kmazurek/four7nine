magic
tech scmos
timestamp 1385337736
<< pwell >>
rect -150 -113 -94 -99
rect -149 -125 -94 -113
rect -150 -197 -94 -175
rect -26 -197 8 -179
<< nwell >>
rect -150 -89 -94 -57
rect -150 -165 -94 -143
rect -26 -157 -3 -143
<< polysilicon >>
rect -120 -76 -116 -74
rect -106 -76 -102 -74
rect -142 -84 -138 -82
rect -142 -92 -138 -88
rect -142 -100 -138 -96
rect -120 -100 -116 -80
rect -142 -106 -138 -104
rect -120 -108 -116 -104
rect -106 -87 -102 -80
rect -106 -108 -102 -91
rect -94 -104 -83 -100
rect -120 -114 -116 -112
rect -106 -114 -102 -112
rect -95 -124 -63 -120
rect -120 -152 -116 -150
rect -106 -152 -102 -150
rect -18 -152 -14 -150
rect -142 -160 -138 -158
rect -142 -168 -138 -164
rect -142 -176 -138 -172
rect -120 -176 -116 -156
rect -142 -182 -138 -180
rect -120 -184 -116 -180
rect -106 -163 -102 -156
rect -106 -184 -102 -167
rect -18 -168 -14 -156
rect -18 -184 -14 -172
rect -120 -190 -116 -188
rect -106 -190 -102 -188
rect -18 -190 -14 -188
<< ndiffusion >>
rect -145 -104 -142 -100
rect -138 -104 -135 -100
rect -123 -112 -120 -108
rect -116 -112 -106 -108
rect -102 -112 -99 -108
rect -145 -180 -142 -176
rect -138 -180 -135 -176
rect -123 -188 -120 -184
rect -116 -188 -106 -184
rect -102 -188 -99 -184
rect -21 -188 -18 -184
rect -14 -188 -11 -184
<< pdiffusion >>
rect -123 -80 -120 -76
rect -116 -80 -113 -76
rect -109 -80 -106 -76
rect -102 -80 -99 -76
rect -145 -88 -142 -84
rect -138 -88 -135 -84
rect -123 -156 -120 -152
rect -116 -156 -113 -152
rect -109 -156 -106 -152
rect -102 -156 -99 -152
rect -21 -156 -18 -152
rect -14 -156 -11 -152
rect -145 -164 -142 -160
rect -138 -164 -135 -160
<< metal1 >>
rect -21 -47 110 -43
rect -21 -50 -17 -47
rect 5 -54 69 -50
rect -150 -62 -149 -58
rect -136 -62 -90 -58
rect -86 -62 -63 -58
rect -135 -84 -131 -62
rect -127 -76 -123 -62
rect -99 -76 -95 -62
rect 65 -78 69 -54
rect -149 -92 -145 -88
rect -113 -92 -109 -80
rect -102 -91 -86 -87
rect -157 -96 -145 -92
rect -138 -96 -109 -92
rect -149 -100 -145 -96
rect -135 -120 -131 -104
rect -127 -108 -123 -96
rect -116 -104 -98 -100
rect -99 -120 -95 -112
rect -150 -124 -149 -120
rect -136 -124 -99 -120
rect -90 -128 -86 -91
rect -79 -104 -75 -100
rect 65 -128 69 -82
rect 106 -102 110 -47
rect 106 -106 114 -102
rect 106 -128 110 -106
rect -90 -132 65 -128
rect 91 -132 110 -128
rect -157 -140 -47 -136
rect -3 -140 23 -136
rect -3 -144 1 -140
rect -150 -148 -149 -144
rect -136 -148 -90 -144
rect -86 -148 -15 -144
rect -4 -148 1 -144
rect -135 -160 -131 -148
rect -127 -152 -123 -148
rect -99 -152 -95 -148
rect -11 -152 -7 -148
rect -149 -168 -145 -164
rect -113 -168 -109 -156
rect -102 -167 -75 -163
rect -25 -168 -21 -156
rect -157 -172 -145 -168
rect -138 -172 -109 -168
rect -43 -172 -21 -168
rect -14 -172 14 -168
rect -149 -176 -145 -172
rect -135 -192 -131 -180
rect -127 -184 -123 -172
rect -116 -180 -112 -176
rect -99 -192 -95 -188
rect -150 -196 -149 -192
rect -136 -196 -94 -192
rect -81 -206 -77 -180
rect -25 -184 -21 -172
rect 10 -182 14 -172
rect -11 -192 -7 -188
rect -69 -196 -55 -192
rect -51 -196 -25 -192
rect -14 -196 12 -192
rect 8 -198 12 -196
rect 8 -202 23 -198
rect 106 -206 110 -132
rect -81 -210 110 -206
<< metal2 >>
rect -90 -144 -86 -62
rect 69 -82 114 -78
rect -75 -163 -71 -104
rect -108 -180 -81 -176
rect -55 -192 -51 -124
rect -47 -168 -43 -140
rect -90 -196 -73 -192
<< ntransistor >>
rect -142 -104 -138 -100
rect -120 -112 -116 -108
rect -106 -112 -102 -108
rect -142 -180 -138 -176
rect -120 -188 -116 -184
rect -106 -188 -102 -184
rect -18 -188 -14 -184
<< ptransistor >>
rect -120 -80 -116 -76
rect -106 -80 -102 -76
rect -142 -88 -138 -84
rect -120 -156 -116 -152
rect -106 -156 -102 -152
rect -18 -156 -14 -152
rect -142 -164 -138 -160
<< polycontact >>
rect -21 -54 -17 -50
rect 1 -54 5 -50
rect -142 -96 -138 -92
rect -120 -104 -116 -100
rect -106 -91 -102 -87
rect -98 -104 -94 -100
rect -83 -104 -79 -100
rect -99 -124 -95 -120
rect -63 -124 -59 -120
rect 65 -132 69 -128
rect 87 -132 91 -128
rect -142 -172 -138 -168
rect -120 -180 -116 -176
rect -106 -167 -102 -163
rect -18 -172 -14 -168
<< ndcontact >>
rect -149 -104 -145 -100
rect -135 -104 -131 -100
rect -127 -112 -123 -108
rect -99 -112 -95 -108
rect -149 -180 -145 -176
rect -135 -180 -131 -176
rect -127 -188 -123 -184
rect -99 -188 -95 -184
rect -25 -188 -21 -184
rect -11 -188 -7 -184
<< pdcontact >>
rect -127 -80 -123 -76
rect -113 -80 -109 -76
rect -99 -80 -95 -76
rect -149 -88 -145 -84
rect -135 -88 -131 -84
rect -127 -156 -123 -152
rect -113 -156 -109 -152
rect -99 -156 -95 -152
rect -25 -156 -21 -152
rect -11 -156 -7 -152
rect -149 -164 -145 -160
rect -135 -164 -131 -160
<< m2contact >>
rect -90 -62 -86 -58
rect 65 -82 69 -78
rect -75 -104 -71 -100
rect -55 -124 -51 -120
rect -47 -140 -43 -136
rect -90 -148 -86 -144
rect -75 -167 -71 -163
rect -47 -172 -43 -168
rect -112 -180 -108 -176
rect -81 -180 -77 -176
rect -94 -196 -90 -192
rect -73 -196 -69 -192
rect -55 -196 -51 -192
<< psubstratepcontact >>
rect -149 -124 -136 -120
rect -149 -196 -136 -192
rect -25 -196 -14 -192
<< nsubstratencontact >>
rect -149 -62 -136 -58
rect -149 -148 -136 -144
rect -15 -148 -4 -144
use XOR  XOR_0
timestamp 1385331530
transform -1 0 -4 0 1 -78
box -20 -47 68 24
use XOR  XOR_1
timestamp 1385331530
transform -1 0 82 0 1 -156
box -20 -47 68 24
<< labels >>
rlabel metal1 -156 -138 -156 -138 3 Out00
rlabel metal1 -82 -59 -82 -59 5 Vdd
rlabel metal1 -83 -145 -83 -145 5 Vdd
rlabel metal1 -65 -195 -65 -195 1 GND
rlabel metal1 -156 -94 -156 -94 3 Out10
rlabel metal1 -156 -170 -156 -170 3 Out01
rlabel metal2 113 -80 113 -80 7 Sel0
rlabel metal1 113 -104 113 -104 7 Sel1
<< end >>
