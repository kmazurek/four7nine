magic
tech scmos
timestamp 1385158978
<< pwell >>
rect 4 -17 46 3
rect -60 -43 46 -17
<< nwell >>
rect -60 -5 -18 27
<< polysilicon >>
rect 5 10 9 30
rect 23 2 27 30
rect -52 0 -48 2
rect -30 0 -26 2
rect -52 -8 -48 -4
rect -52 -16 -48 -12
rect -30 -8 -26 -4
rect 1 -9 5 -5
rect 9 -9 11 -5
rect 41 -6 45 30
rect -30 -16 -26 -12
rect 19 -17 23 -13
rect 27 -17 29 -13
rect -52 -22 -48 -20
rect -30 -22 -26 -20
rect 37 -25 41 -21
rect 45 -25 47 -21
<< ndiffusion >>
rect 5 -5 9 -2
rect 5 -12 9 -9
rect 23 -13 27 -10
rect -55 -20 -52 -16
rect -48 -20 -45 -16
rect -33 -20 -30 -16
rect -26 -20 -23 -16
rect 23 -20 27 -17
rect 41 -21 45 -18
rect 41 -28 45 -25
<< pdiffusion >>
rect -55 -4 -52 0
rect -48 -4 -45 0
rect -33 -4 -30 0
rect -26 -4 -23 0
<< metal1 >>
rect -62 22 -59 26
rect -46 22 49 26
rect -45 0 -41 22
rect -23 0 -19 22
rect -3 14 53 18
rect -59 -8 -55 -4
rect -37 -8 -33 -4
rect -3 -5 1 14
rect 5 2 9 6
rect 15 6 53 10
rect -63 -12 -55 -8
rect -48 -12 -33 -8
rect -26 -12 -11 -8
rect -59 -16 -55 -12
rect -37 -16 -33 -12
rect -15 -16 5 -12
rect 15 -13 19 6
rect 23 -6 27 -2
rect 33 -2 53 2
rect -45 -38 -41 -20
rect -23 -38 -19 -20
rect -15 -20 -11 -16
rect -15 -24 23 -20
rect 33 -21 37 -2
rect 41 -14 45 -10
rect -15 -28 -11 -24
rect -15 -32 41 -28
rect -62 -42 -59 -38
rect -46 -42 51 -38
<< ntransistor >>
rect 5 -9 9 -5
rect -52 -20 -48 -16
rect -30 -20 -26 -16
rect 23 -17 27 -13
rect 41 -25 45 -21
<< ptransistor >>
rect -52 -4 -48 0
rect -30 -4 -26 0
<< polycontact >>
rect 5 6 9 10
rect 23 -2 27 2
rect -52 -12 -48 -8
rect -30 -12 -26 -8
rect -3 -9 1 -5
rect 41 -10 45 -6
rect 15 -17 19 -13
rect 33 -25 37 -21
<< ndcontact >>
rect 5 -2 9 2
rect 5 -16 9 -12
rect 23 -10 27 -6
rect -59 -20 -55 -16
rect -45 -20 -41 -16
rect -37 -20 -33 -16
rect -23 -20 -19 -16
rect 23 -24 27 -20
rect 41 -18 45 -14
rect 41 -32 45 -28
<< pdcontact >>
rect -59 -4 -55 0
rect -45 -4 -41 0
rect -37 -4 -33 0
rect -23 -4 -19 0
<< psubstratepcontact >>
rect -59 -42 -46 -38
<< nsubstratencontact >>
rect -59 22 -46 26
<< labels >>
rlabel metal1 -21 25 -21 25 5 Vdd
rlabel metal1 -62 -10 -62 -10 3 Out
rlabel metal1 -21 -41 -21 -41 1 GND
rlabel metal1 52 16 52 16 7 Sel0
rlabel metal1 52 8 52 8 7 Sel1
rlabel metal1 52 0 52 0 7 Sel2
rlabel polysilicon 7 29 7 29 5 In0
rlabel polysilicon 25 29 25 29 5 In1
rlabel polysilicon 43 29 43 29 5 In2
<< end >>
