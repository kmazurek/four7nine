magic
tech scmos
timestamp 1386045209
<< polysilicon >>
rect -36 -131 129 -129
<< metal1 >>
rect -36 165 9 169
rect -37 156 8 160
rect -34 148 135 152
rect -16 22 119 26
rect 351 -8 396 -4
rect 351 -16 396 -12
rect 352 -24 397 -20
rect -34 -66 129 -59
<< metal2 >>
rect 345 -76 390 -72
rect 351 -104 396 -100
rect 300 -139 396 -135
use mux1  mux1_0
timestamp 1385976061
transform 1 0 127 0 1 6
box -127 -110 275 678
use shift1  shift1_0
timestamp 1385976061
transform 1 0 -35 0 1 -163
box -3 12 417 315
use reg1  reg1_0
timestamp 1386043477
transform 1 0 62 0 1 -365
box -82 213 332 474
<< labels >>
rlabel metal1 -37 156 8 160 1 sel0
rlabel metal1 351 -8 396 -4 1 inbit
rlabel metal1 351 -16 396 -12 1 inbit_next
rlabel metal1 352 -24 397 -20 1 shift
rlabel metal2 345 -76 390 -72 1 clk
rlabel metal2 351 -104 396 -100 1 Qout1
rlabel space 298 -139 394 -135 3 rst
rlabel metal2 300 -139 396 -135 3 rst
rlabel polysilicon -36 -131 129 -129 7 Din
rlabel metal1 -36 165 9 169 1 sel1
rlabel metal1 -34 148 135 152 5 Vdd
rlabel space -16 -151 130 -144 7 GND
rlabel space 20 86 119 90 1 Vdd
rlabel space 31 18 105 25 1 GND
rlabel metal1 -34 -66 129 -59 5 Vd
<< end >>
