magic
tech scmos
timestamp 1385338104
<< polysilicon >>
rect -56 88 -52 92
rect -38 88 -34 92
rect -20 88 -16 92
<< metal1 >>
rect -8 142 7 146
rect -4 76 0 112
rect 271 98 275 102
rect -14 72 0 76
rect -14 64 0 68
rect -14 56 0 60
rect -128 46 -124 50
rect -4 32 0 56
rect -12 12 -8 20
rect -12 8 7 12
<< metal2 >>
rect -12 84 -8 142
rect 271 122 275 126
<< m2contact >>
rect -12 142 -8 146
rect -12 80 -8 84
use 31MUX  31MUX_0
timestamp 1385158978
transform 1 0 -61 0 1 58
box -63 -43 53 30
use MUXsel  MUXsel_0
timestamp 1385337736
transform 1 0 157 0 1 204
box -157 -210 114 -43
<< labels >>
rlabel metal1 -1 145 -1 145 5 Vdd
rlabel metal1 -5 9 -5 9 1 GND
rlabel polysilicon -54 91 -54 91 5 In0
rlabel polysilicon -36 91 -36 91 5 In1
rlabel polysilicon -18 91 -18 91 5 In2
rlabel metal1 -127 48 -127 48 3 Out
rlabel metal2 274 124 274 124 7 Sel0
rlabel metal1 274 100 274 100 7 Sel1
<< end >>
