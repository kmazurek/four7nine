magic
tech scmos
timestamp 1385600620
<< pwell >>
rect 56 91 299 127
<< nwell >>
rect 56 127 299 178
<< polysilicon >>
rect 70 137 72 152
rect 87 137 89 161
rect 103 137 105 152
rect 121 137 123 139
rect 131 137 133 173
rect 189 140 191 156
rect 149 137 151 139
rect 169 138 191 140
rect 169 137 171 138
rect 189 137 191 138
rect 211 137 213 139
rect 236 137 238 139
rect 260 137 262 139
rect 270 137 272 173
rect 286 137 288 156
rect 70 120 72 133
rect 87 120 89 133
rect 103 131 105 133
rect 103 120 105 122
rect 121 120 123 133
rect 131 120 133 133
rect 149 120 151 133
rect 169 130 171 133
rect 189 128 191 133
rect 169 120 171 123
rect 189 120 191 122
rect 211 120 213 133
rect 236 120 238 133
rect 260 120 262 133
rect 270 120 272 133
rect 286 131 288 133
rect 286 120 288 123
rect 70 114 72 116
rect 87 114 89 116
rect 103 92 105 116
rect 121 114 123 116
rect 131 114 133 116
rect 149 114 151 116
rect 169 115 171 116
rect 189 115 191 116
rect 169 113 191 115
rect 211 114 213 116
rect 236 114 238 116
rect 169 92 171 113
rect 260 111 262 116
rect 270 114 272 116
rect 252 107 262 111
rect 286 92 288 116
<< ndiffusion >>
rect 69 116 70 120
rect 72 116 73 120
rect 86 116 87 120
rect 89 116 90 120
rect 102 116 103 120
rect 105 116 106 120
rect 120 116 121 120
rect 123 116 125 120
rect 129 116 131 120
rect 133 116 134 120
rect 148 116 149 120
rect 151 116 152 120
rect 168 116 169 120
rect 171 116 172 120
rect 188 116 189 120
rect 191 116 192 120
rect 210 116 211 120
rect 213 116 214 120
rect 235 116 236 120
rect 238 116 239 120
rect 259 116 260 120
rect 262 116 264 120
rect 268 116 270 120
rect 272 116 273 120
rect 285 116 286 120
rect 288 116 289 120
<< pdiffusion >>
rect 69 133 70 137
rect 72 133 73 137
rect 86 133 87 137
rect 89 133 90 137
rect 102 133 103 137
rect 105 133 106 137
rect 120 133 121 137
rect 123 133 131 137
rect 133 133 134 137
rect 148 133 149 137
rect 151 133 152 137
rect 168 133 169 137
rect 171 133 172 137
rect 188 133 189 137
rect 191 133 192 137
rect 210 133 211 137
rect 213 133 214 137
rect 235 133 236 137
rect 238 133 239 137
rect 259 133 260 137
rect 262 133 270 137
rect 272 133 273 137
rect 285 133 286 137
rect 288 133 289 137
<< metal1 >>
rect 133 173 266 177
rect 272 173 298 177
rect 57 161 83 165
rect 76 152 102 156
rect 114 152 191 156
rect 199 152 288 156
rect 86 141 201 145
rect 260 141 298 145
rect 73 140 298 141
rect 73 137 77 140
rect 82 137 86 140
rect 116 137 120 140
rect 144 137 148 140
rect 206 137 210 140
rect 231 137 235 140
rect 255 137 259 140
rect 65 120 69 133
rect 90 127 94 133
rect 98 127 102 133
rect 90 123 102 127
rect 90 120 94 123
rect 73 104 77 116
rect 98 120 102 123
rect 106 130 110 133
rect 110 126 117 130
rect 134 127 138 133
rect 152 127 156 133
rect 164 127 168 133
rect 106 120 110 126
rect 125 123 139 127
rect 143 123 145 127
rect 152 123 168 127
rect 125 120 129 123
rect 152 120 156 123
rect 82 104 86 116
rect 116 104 120 116
rect 134 104 138 116
rect 164 120 168 123
rect 172 127 176 133
rect 172 120 176 123
rect 184 127 188 133
rect 184 120 188 123
rect 192 127 196 133
rect 214 127 218 133
rect 239 127 243 133
rect 246 127 250 131
rect 273 127 277 133
rect 281 127 285 133
rect 192 123 200 127
rect 204 123 207 127
rect 214 123 232 127
rect 239 123 250 127
rect 264 123 285 127
rect 289 127 293 133
rect 192 120 196 123
rect 214 120 218 123
rect 144 104 148 116
rect 206 104 210 116
rect 222 111 226 123
rect 239 120 243 123
rect 264 120 268 123
rect 281 120 285 123
rect 231 104 235 116
rect 243 107 248 111
rect 255 104 259 116
rect 273 104 277 116
rect 95 100 107 104
rect 154 100 222 104
rect 262 100 298 104
rect 57 92 61 96
rect 65 92 95 96
rect 103 92 165 96
rect 169 92 282 96
rect 286 92 298 96
<< metal2 >>
rect 246 159 298 163
rect 106 147 176 151
rect 106 130 110 147
rect 172 127 176 147
rect 246 135 250 159
rect 61 96 65 122
rect 139 112 143 123
rect 180 112 184 127
rect 192 116 196 120
rect 139 108 184 112
rect 200 100 204 123
rect 226 107 239 111
rect 289 100 293 123
rect 200 96 293 100
<< ntransistor >>
rect 70 116 72 120
rect 87 116 89 120
rect 103 116 105 120
rect 121 116 123 120
rect 131 116 133 120
rect 149 116 151 120
rect 169 116 171 120
rect 189 116 191 120
rect 211 116 213 120
rect 236 116 238 120
rect 260 116 262 120
rect 270 116 272 120
rect 286 116 288 120
<< ptransistor >>
rect 70 133 72 137
rect 87 133 89 137
rect 103 133 105 137
rect 121 133 123 137
rect 131 133 133 137
rect 149 133 151 137
rect 169 133 171 137
rect 189 133 191 137
rect 211 133 213 137
rect 236 133 238 137
rect 260 133 262 137
rect 270 133 272 137
rect 286 133 288 137
<< polycontact >>
rect 123 173 133 177
rect 266 173 272 177
rect 83 161 89 165
rect 70 152 76 156
rect 102 152 114 156
rect 191 152 199 156
rect 288 152 294 156
rect 117 126 121 130
rect 145 123 149 127
rect 207 123 211 127
rect 232 123 236 127
rect 95 92 103 96
rect 165 92 169 96
rect 248 107 252 111
rect 282 92 286 96
<< ndcontact >>
rect 65 116 69 120
rect 73 116 77 120
rect 82 116 86 120
rect 90 116 94 120
rect 98 116 102 120
rect 106 116 110 120
rect 116 116 120 120
rect 125 116 129 120
rect 134 116 138 120
rect 144 116 148 120
rect 152 116 156 120
rect 164 116 168 120
rect 172 116 176 120
rect 184 116 188 120
rect 192 116 196 120
rect 206 116 210 120
rect 214 116 218 120
rect 231 116 235 120
rect 239 116 243 120
rect 255 116 259 120
rect 264 116 268 120
rect 273 116 277 120
rect 281 116 285 120
rect 289 116 293 120
<< pdcontact >>
rect 65 133 69 137
rect 73 133 77 137
rect 82 133 86 137
rect 90 133 94 137
rect 98 133 102 137
rect 106 133 110 137
rect 116 133 120 137
rect 134 133 138 137
rect 144 133 148 137
rect 152 133 156 137
rect 164 133 168 137
rect 172 133 176 137
rect 184 133 188 137
rect 192 133 196 137
rect 206 133 210 137
rect 214 133 218 137
rect 231 133 235 137
rect 239 133 243 137
rect 255 133 259 137
rect 273 133 277 137
rect 281 133 285 137
rect 289 133 293 137
<< m2contact >>
rect 61 122 65 126
rect 106 126 110 130
rect 139 123 143 127
rect 172 123 176 127
rect 184 123 188 127
rect 246 131 250 135
rect 200 123 204 127
rect 289 123 293 127
rect 222 107 226 111
rect 239 107 243 111
rect 61 92 65 96
<< psubstratepcontact >>
rect 73 100 95 104
rect 107 100 154 104
rect 222 100 262 104
<< nsubstratencontact >>
rect 73 141 86 145
rect 201 141 260 145
<< labels >>
rlabel metal1 57 94 57 94 7 clkb
rlabel metal1 98 101 98 101 1 GND
rlabel metal1 95 144 95 144 5 Vdd
rlabel metal1 279 155 279 155 5 clk
rlabel metal1 57 163 57 163 7 D
rlabel metal1 298 175 298 175 3 rst
rlabel metal2 298 161 298 161 3 Q
<< end >>
