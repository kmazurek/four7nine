magic
tech scmos
timestamp 1386052290
<< pwell >>
rect 30 132 281 186
rect 175 88 227 92
rect 93 48 227 88
rect 38 -71 66 -61
rect 76 -90 246 -76
rect 76 -95 261 -90
rect 46 -114 261 -95
rect 175 -446 257 -436
rect 94 -464 150 -450
rect 95 -476 150 -464
rect 200 -476 257 -446
rect 30 -514 72 -494
rect -29 -540 72 -514
rect 229 -523 311 -514
rect 94 -548 150 -526
rect 227 -530 311 -523
rect 186 -548 311 -530
rect 187 -554 311 -548
rect -41 -594 90 -561
rect 56 -752 307 -698
<< nwell >>
rect 31 193 282 247
rect 93 102 227 116
rect 93 98 185 102
rect 38 -53 246 -33
rect 76 -66 246 -53
rect 35 -87 66 -77
rect 94 -440 150 -408
rect 215 -426 257 -408
rect -29 -502 13 -470
rect 94 -516 150 -494
rect 186 -508 209 -494
rect 269 -504 311 -486
rect -41 -637 90 -594
rect -41 -638 308 -637
rect 57 -691 308 -638
<< polysilicon >>
rect -12 53 -7 239
rect 7 165 9 268
rect 46 210 77 212
rect 46 203 48 210
rect 69 203 71 207
rect 81 203 83 212
rect 90 205 105 207
rect 103 203 105 205
rect 114 203 116 206
rect 137 203 139 205
rect 189 203 191 210
rect 216 203 218 205
rect 227 203 229 205
rect 240 203 242 205
rect 267 203 269 206
rect 46 177 48 195
rect 46 175 51 177
rect 55 175 57 177
rect 69 165 71 195
rect 81 192 83 195
rect 103 174 105 195
rect 114 174 116 195
rect 137 187 139 195
rect 124 185 139 187
rect 137 173 139 185
rect 151 180 153 189
rect 177 185 179 193
rect 177 178 179 181
rect 151 173 153 176
rect 137 171 142 173
rect 146 171 148 173
rect 189 173 191 195
rect 216 185 218 195
rect 198 183 218 185
rect 216 174 218 183
rect 227 174 229 195
rect 240 185 242 195
rect 186 171 194 173
rect 198 171 200 173
rect 103 167 105 170
rect 7 163 74 165
rect 78 163 80 165
rect 114 163 116 170
rect 267 173 269 195
rect 249 171 272 173
rect 276 171 280 173
rect 216 167 218 170
rect 227 163 229 170
rect 101 107 105 123
rect 127 119 256 123
rect 123 103 127 119
rect 193 107 197 109
rect 215 107 219 109
rect 256 104 260 119
rect 101 95 105 103
rect 193 99 197 103
rect 101 87 105 91
rect 101 71 105 83
rect 123 79 127 99
rect 193 91 197 95
rect 215 99 219 103
rect 215 91 219 95
rect 123 63 127 75
rect 146 63 150 91
rect 163 87 167 89
rect 193 85 197 87
rect 215 85 219 87
rect 163 71 167 83
rect 146 57 150 59
rect 162 -19 166 41
rect 46 -45 50 -43
rect 84 -44 88 -23
rect 91 -44 95 -31
rect 98 -44 102 -42
rect 120 -44 124 -42
rect 148 -44 152 -31
rect 162 -44 166 -23
rect 196 -44 200 -31
rect 203 -44 207 -23
rect 235 -27 239 95
rect 235 -44 239 -31
rect 249 -44 253 -23
rect 46 -56 50 -49
rect 46 -64 50 -60
rect 46 -70 50 -68
rect 54 -80 58 -78
rect 54 -88 58 -84
rect 84 -91 88 -48
rect 91 -91 95 -48
rect 98 -61 102 -48
rect 98 -91 102 -65
rect 120 -61 124 -48
rect 134 -61 138 -59
rect 120 -91 124 -65
rect 134 -69 138 -65
rect 134 -77 138 -73
rect 134 -83 138 -81
rect 54 -96 58 -92
rect 148 -95 152 -48
rect 162 -95 166 -48
rect 196 -91 200 -48
rect 203 -91 207 -48
rect 221 -55 225 -53
rect 221 -69 225 -59
rect 221 -83 225 -73
rect 221 -89 225 -87
rect 235 -91 239 -48
rect 249 -91 253 -48
rect 84 -97 88 -95
rect 91 -97 95 -95
rect 98 -97 102 -95
rect 120 -97 124 -95
rect 196 -97 200 -95
rect 203 -97 207 -95
rect 235 -97 239 -95
rect 249 -97 253 -95
rect 54 -102 58 -100
rect 148 -103 152 -99
rect 162 -103 166 -99
rect 31 -487 35 -139
rect 49 -495 53 -130
rect -21 -497 -17 -495
rect 1 -497 5 -495
rect 67 -143 71 -135
rect -21 -505 -17 -501
rect -21 -513 -17 -509
rect 1 -505 5 -501
rect 27 -506 31 -502
rect 35 -506 37 -502
rect 67 -503 71 -147
rect 223 -421 227 -405
rect 245 -417 249 -405
rect 124 -427 128 -425
rect 138 -427 142 -425
rect 102 -435 106 -433
rect 102 -443 106 -439
rect 102 -451 106 -447
rect 124 -451 128 -431
rect 102 -457 106 -455
rect 124 -459 128 -455
rect 138 -438 142 -431
rect 183 -437 187 -435
rect 138 -459 142 -442
rect 150 -455 161 -451
rect 183 -453 187 -441
rect 200 -461 204 -433
rect 223 -445 227 -425
rect 245 -437 249 -421
rect 223 -461 227 -449
rect 245 -453 249 -441
rect 124 -465 128 -463
rect 138 -465 142 -463
rect 200 -467 204 -465
rect 149 -475 181 -471
rect 277 -499 281 -483
rect 299 -495 303 -483
rect 124 -503 128 -501
rect 138 -503 142 -501
rect 194 -503 198 -501
rect 1 -513 5 -509
rect 45 -514 49 -510
rect 53 -514 55 -510
rect 102 -511 106 -509
rect -21 -519 -17 -517
rect 1 -519 5 -517
rect 63 -522 67 -518
rect 71 -522 73 -518
rect 102 -519 106 -515
rect 102 -527 106 -523
rect 124 -527 128 -507
rect 102 -533 106 -531
rect 124 -535 128 -531
rect 138 -514 142 -507
rect 138 -535 142 -518
rect 194 -519 198 -507
rect 237 -515 241 -513
rect 194 -535 198 -523
rect 237 -531 241 -519
rect 254 -539 258 -511
rect 277 -523 281 -503
rect 299 -515 303 -499
rect 277 -539 281 -527
rect 124 -541 128 -539
rect 138 -541 142 -539
rect 194 -541 198 -539
rect 299 -531 303 -519
rect 254 -545 258 -543
rect 299 -557 303 -535
rect 69 -576 71 -574
rect 39 -578 51 -576
rect -22 -584 -20 -582
rect -2 -584 0 -582
rect 18 -584 20 -582
rect 39 -584 41 -578
rect 58 -584 60 -582
rect -22 -604 -20 -588
rect -22 -620 -20 -608
rect -2 -613 0 -588
rect 18 -595 20 -588
rect -2 -620 0 -617
rect 18 -620 20 -599
rect 39 -620 41 -588
rect 58 -603 60 -588
rect 69 -603 71 -580
rect 58 -609 60 -607
rect 69 -620 71 -607
rect -22 -626 -20 -624
rect -2 -626 0 -624
rect 18 -626 20 -624
rect 39 -626 41 -624
rect 69 -626 71 -624
rect 72 -674 103 -672
rect 72 -681 74 -674
rect 95 -681 97 -677
rect 107 -681 109 -672
rect 116 -679 131 -677
rect 129 -681 131 -679
rect 140 -681 142 -678
rect 163 -681 165 -679
rect 215 -681 217 -674
rect 242 -681 244 -679
rect 253 -681 255 -679
rect 266 -681 268 -679
rect 293 -681 295 -678
rect 72 -707 74 -689
rect 72 -709 77 -707
rect 81 -709 83 -707
rect 95 -719 97 -689
rect 107 -692 109 -689
rect 129 -710 131 -689
rect 140 -710 142 -689
rect 163 -697 165 -689
rect 150 -699 165 -697
rect 163 -711 165 -699
rect 177 -704 179 -695
rect 203 -699 205 -691
rect 203 -706 205 -703
rect 177 -711 179 -708
rect 163 -713 168 -711
rect 172 -713 174 -711
rect 215 -711 217 -689
rect 242 -699 244 -689
rect 224 -701 244 -699
rect 242 -710 244 -701
rect 253 -710 255 -689
rect 266 -699 268 -689
rect 212 -713 220 -711
rect 224 -713 226 -711
rect 129 -717 131 -714
rect 42 -721 100 -719
rect 104 -721 106 -719
rect 140 -721 142 -714
rect 293 -711 295 -689
rect 275 -713 298 -711
rect 302 -713 306 -711
rect 242 -717 244 -714
rect 253 -721 255 -714
<< ndiffusion >>
rect 51 177 55 180
rect 51 172 55 175
rect 100 170 103 174
rect 105 170 107 174
rect 111 170 114 174
rect 116 170 120 174
rect 174 181 177 185
rect 179 181 182 185
rect 146 176 151 180
rect 153 176 156 180
rect 142 173 146 176
rect 194 173 198 176
rect 74 165 78 168
rect 142 168 146 171
rect 194 168 198 171
rect 213 170 216 174
rect 218 170 220 174
rect 224 170 227 174
rect 229 170 233 174
rect 272 173 276 176
rect 272 168 276 171
rect 74 160 78 163
rect 98 83 101 87
rect 105 83 108 87
rect 120 75 123 79
rect 127 75 130 79
rect 190 87 193 91
rect 197 87 200 91
rect 212 87 215 91
rect 219 87 222 91
rect 160 83 163 87
rect 167 83 170 87
rect 143 59 146 63
rect 150 59 153 63
rect 43 -68 46 -64
rect 50 -68 53 -64
rect 131 -81 134 -77
rect 138 -81 141 -77
rect 81 -95 84 -91
rect 88 -95 91 -91
rect 95 -95 98 -91
rect 102 -95 105 -91
rect 117 -95 120 -91
rect 124 -95 127 -91
rect 218 -87 221 -83
rect 225 -87 228 -83
rect 193 -95 196 -91
rect 200 -95 203 -91
rect 207 -95 210 -91
rect 232 -95 235 -91
rect 239 -95 242 -91
rect 246 -95 249 -91
rect 253 -95 256 -91
rect 51 -100 54 -96
rect 58 -100 61 -96
rect 144 -99 148 -95
rect 152 -99 155 -95
rect 159 -99 162 -95
rect 166 -99 169 -95
rect 31 -502 35 -499
rect 99 -455 102 -451
rect 106 -455 109 -451
rect 180 -441 183 -437
rect 187 -441 190 -437
rect 121 -463 124 -459
rect 128 -463 138 -459
rect 142 -463 145 -459
rect 242 -441 245 -437
rect 249 -441 252 -437
rect 220 -449 223 -445
rect 227 -449 230 -445
rect 197 -465 200 -461
rect 204 -465 207 -461
rect 31 -509 35 -506
rect 49 -510 53 -507
rect -24 -517 -21 -513
rect -17 -517 -14 -513
rect -2 -517 1 -513
rect 5 -517 8 -513
rect 49 -517 53 -514
rect 67 -518 71 -515
rect 67 -525 71 -522
rect 99 -531 102 -527
rect 106 -531 109 -527
rect 234 -519 237 -515
rect 241 -519 244 -515
rect 121 -539 124 -535
rect 128 -539 138 -535
rect 142 -539 145 -535
rect 191 -539 194 -535
rect 198 -539 201 -535
rect 296 -519 299 -515
rect 303 -519 306 -515
rect 274 -527 277 -523
rect 281 -527 284 -523
rect 251 -543 254 -539
rect 258 -543 261 -539
rect 67 -580 69 -576
rect 71 -580 73 -576
rect -25 -588 -22 -584
rect -20 -588 -17 -584
rect -5 -588 -2 -584
rect 0 -588 3 -584
rect 15 -588 18 -584
rect 20 -588 23 -584
rect 36 -588 39 -584
rect 41 -588 44 -584
rect 56 -588 58 -584
rect 60 -588 62 -584
rect 77 -707 81 -704
rect 77 -712 81 -709
rect 126 -714 129 -710
rect 131 -714 133 -710
rect 137 -714 140 -710
rect 142 -714 146 -710
rect 200 -703 203 -699
rect 205 -703 208 -699
rect 172 -708 177 -704
rect 179 -708 182 -704
rect 168 -711 172 -708
rect 220 -711 224 -708
rect 100 -719 104 -716
rect 168 -716 172 -713
rect 220 -716 224 -713
rect 239 -714 242 -710
rect 244 -714 246 -710
rect 250 -714 253 -710
rect 255 -714 259 -710
rect 298 -711 302 -708
rect 298 -716 302 -713
rect 100 -724 104 -721
<< pdiffusion >>
rect 43 195 46 203
rect 48 195 51 203
rect 66 195 69 203
rect 71 195 74 203
rect 78 195 81 203
rect 83 195 86 203
rect 100 195 103 203
rect 105 195 114 203
rect 116 195 120 203
rect 134 195 137 203
rect 139 195 142 203
rect 186 195 189 203
rect 191 195 194 203
rect 213 195 216 203
rect 218 195 227 203
rect 229 195 233 203
rect 237 195 240 203
rect 242 195 245 203
rect 264 195 267 203
rect 269 195 272 203
rect 98 103 101 107
rect 105 103 108 107
rect 190 103 193 107
rect 197 103 200 107
rect 212 103 215 107
rect 219 103 222 107
rect 120 99 123 103
rect 127 99 130 103
rect 43 -49 46 -45
rect 50 -49 53 -45
rect 81 -48 84 -44
rect 88 -48 91 -44
rect 95 -48 98 -44
rect 102 -48 105 -44
rect 117 -48 120 -44
rect 124 -48 128 -44
rect 144 -48 148 -44
rect 152 -48 155 -44
rect 159 -48 162 -44
rect 166 -48 169 -44
rect 193 -48 196 -44
rect 200 -48 203 -44
rect 207 -48 210 -44
rect 232 -48 235 -44
rect 239 -48 242 -44
rect 246 -48 249 -44
rect 253 -48 256 -44
rect 51 -84 54 -80
rect 58 -84 61 -80
rect 131 -65 134 -61
rect 138 -65 141 -61
rect 218 -59 221 -55
rect 225 -59 228 -55
rect -24 -501 -21 -497
rect -17 -501 -14 -497
rect -2 -501 1 -497
rect 5 -501 8 -497
rect 242 -421 245 -417
rect 249 -421 252 -417
rect 220 -425 223 -421
rect 227 -425 230 -421
rect 121 -431 124 -427
rect 128 -431 131 -427
rect 135 -431 138 -427
rect 142 -431 145 -427
rect 99 -439 102 -435
rect 106 -439 109 -435
rect 296 -499 299 -495
rect 303 -499 306 -495
rect 274 -503 277 -499
rect 281 -503 284 -499
rect 121 -507 124 -503
rect 128 -507 131 -503
rect 135 -507 138 -503
rect 142 -507 145 -503
rect 191 -507 194 -503
rect 198 -507 201 -503
rect 99 -515 102 -511
rect 106 -515 109 -511
rect -25 -624 -22 -620
rect -20 -624 -17 -620
rect -5 -624 -2 -620
rect 0 -624 3 -620
rect 15 -624 18 -620
rect 20 -624 23 -620
rect 36 -624 39 -620
rect 41 -624 44 -620
rect 67 -624 69 -620
rect 71 -624 73 -620
rect 69 -689 72 -681
rect 74 -689 77 -681
rect 92 -689 95 -681
rect 97 -689 100 -681
rect 104 -689 107 -681
rect 109 -689 112 -681
rect 126 -689 129 -681
rect 131 -689 140 -681
rect 142 -689 146 -681
rect 160 -689 163 -681
rect 165 -689 168 -681
rect 212 -689 215 -681
rect 217 -689 220 -681
rect 239 -689 242 -681
rect 244 -689 253 -681
rect 255 -689 259 -681
rect 263 -689 266 -681
rect 268 -689 271 -681
rect 290 -689 293 -681
rect 295 -689 298 -681
<< metal1 >>
rect -41 239 -12 247
rect -4 246 321 247
rect -4 239 34 246
rect 270 239 321 246
rect 35 195 39 239
rect 62 203 66 239
rect 77 212 81 218
rect 86 209 90 210
rect 86 203 90 205
rect 96 203 100 239
rect 130 203 134 239
rect 51 184 55 195
rect 39 175 42 179
rect 74 172 78 195
rect 120 181 124 195
rect 107 177 120 181
rect 142 180 146 195
rect 149 193 153 219
rect 107 174 111 177
rect 156 180 160 210
rect 173 193 177 218
rect 182 203 186 239
rect 193 210 194 214
rect 209 203 213 239
rect 245 203 249 206
rect 169 181 170 185
rect 182 175 186 181
rect 194 180 198 195
rect 233 185 237 195
rect 252 189 256 218
rect 260 203 264 239
rect 246 185 256 189
rect 272 188 276 195
rect 220 181 237 185
rect 262 184 276 188
rect 198 176 200 180
rect 220 174 224 181
rect 245 175 249 176
rect 51 136 55 168
rect 74 136 78 156
rect 96 136 100 170
rect 110 159 114 163
rect 120 136 124 170
rect 142 136 146 164
rect 194 136 198 164
rect 209 136 213 170
rect 223 159 227 163
rect 233 136 237 170
rect 262 148 266 184
rect 272 180 276 184
rect 272 136 276 164
rect -41 128 19 136
rect 32 135 322 136
rect 32 128 44 135
rect 280 128 322 135
rect -41 119 123 123
rect 260 119 322 123
rect -41 111 61 115
rect 65 111 109 115
rect 119 111 177 115
rect 181 111 262 115
rect 266 111 322 115
rect 94 107 98 111
rect 108 95 112 103
rect 116 103 120 111
rect 186 107 190 111
rect 208 107 212 111
rect 200 99 204 103
rect 222 99 226 103
rect -41 91 101 95
rect 108 87 112 91
rect 130 87 134 99
rect 178 95 193 99
rect 200 95 215 99
rect 222 95 235 99
rect 142 91 146 95
rect 130 83 156 87
rect 94 53 98 83
rect 130 79 134 83
rect 105 67 109 71
rect 116 53 120 75
rect 170 73 174 83
rect 178 73 182 95
rect 200 91 204 95
rect 222 91 226 95
rect 159 67 163 71
rect 170 69 182 73
rect 170 63 174 69
rect 127 59 139 63
rect 157 59 174 63
rect 186 53 190 87
rect 208 53 212 87
rect 256 78 260 100
rect -41 49 -13 53
rect -5 49 39 53
rect 43 49 98 53
rect 116 49 222 53
rect 226 49 322 53
rect -41 41 162 45
rect 166 41 322 45
rect -41 33 322 37
rect -41 25 322 29
rect -41 17 322 21
rect -41 9 322 13
rect -41 1 322 5
rect -41 -7 322 -3
rect -41 -15 322 -11
rect 88 -23 162 -19
rect 166 -23 203 -19
rect 207 -23 249 -19
rect 61 -35 65 -24
rect 95 -31 148 -27
rect 152 -31 196 -27
rect 200 -31 235 -27
rect -41 -39 117 -35
rect 134 -39 177 -35
rect 181 -39 322 -35
rect 53 -45 57 -39
rect 39 -56 43 -49
rect -40 -60 43 -56
rect 50 -60 53 -56
rect 19 -69 23 -60
rect 39 -64 43 -60
rect 61 -63 65 -39
rect 105 -44 109 -39
rect -41 -73 23 -69
rect 53 -72 57 -68
rect 36 -76 39 -72
rect 43 -76 57 -72
rect 113 -44 117 -39
rect 140 -44 144 -39
rect 169 -44 173 -39
rect 210 -44 214 -39
rect 228 -44 232 -39
rect 256 -44 260 -39
rect 77 -69 81 -48
rect 128 -52 132 -48
rect 128 -56 145 -52
rect 141 -61 145 -56
rect 155 -61 159 -48
rect 102 -65 105 -61
rect 117 -65 120 -61
rect 145 -65 159 -61
rect 127 -69 131 -65
rect 181 -69 185 -64
rect 189 -69 193 -48
rect 242 -55 246 -48
rect 232 -59 246 -55
rect 214 -69 218 -59
rect 36 -79 40 -76
rect 61 -80 65 -69
rect 36 -108 40 -85
rect 69 -73 131 -69
rect 138 -73 218 -69
rect 225 -73 228 -69
rect 232 -73 256 -69
rect 260 -73 322 -69
rect 47 -96 51 -84
rect 69 -88 73 -73
rect 58 -92 73 -88
rect 77 -91 81 -73
rect 127 -77 131 -73
rect 145 -81 159 -77
rect 141 -86 145 -81
rect 127 -90 145 -86
rect 127 -91 131 -90
rect 61 -108 65 -100
rect 105 -108 109 -95
rect 155 -95 159 -81
rect 189 -91 193 -73
rect 214 -83 218 -73
rect 232 -87 246 -83
rect 242 -91 246 -87
rect 113 -108 117 -95
rect 140 -108 144 -99
rect 169 -108 173 -99
rect 210 -108 214 -95
rect 228 -108 232 -95
rect 256 -108 260 -95
rect 36 -112 117 -108
rect 134 -112 241 -108
rect 245 -112 264 -108
rect 268 -112 322 -108
rect 53 -130 159 -126
rect -41 -139 31 -135
rect 35 -139 322 -135
rect -41 -147 67 -143
rect 71 -147 322 -143
rect -41 -155 322 -151
rect -41 -162 322 -158
rect -41 -170 322 -166
rect -41 -178 322 -174
rect -41 -186 322 -182
rect -41 -194 322 -190
rect -41 -202 322 -198
rect -41 -210 322 -206
rect -41 -218 322 -214
rect -41 -226 322 -222
rect -41 -234 322 -230
rect -41 -242 322 -238
rect -41 -250 322 -246
rect -41 -258 322 -254
rect -41 -266 322 -262
rect -41 -274 322 -270
rect -41 -282 322 -278
rect -41 -289 322 -285
rect -41 -297 322 -293
rect -41 -305 322 -301
rect -41 -313 322 -309
rect -41 -321 322 -317
rect -41 -329 322 -325
rect -41 -337 322 -333
rect -41 -345 322 -341
rect -41 -353 322 -349
rect -41 -361 322 -357
rect -41 -369 322 -365
rect -41 -377 322 -373
rect -41 -385 322 -381
rect -41 -396 -29 -392
rect 227 -396 322 -392
rect 223 -401 227 -396
rect -41 -405 -29 -401
rect 249 -405 277 -401
rect -41 -413 -29 -409
rect 79 -413 95 -409
rect 108 -413 154 -409
rect 158 -413 231 -409
rect 241 -413 260 -409
rect 109 -435 113 -413
rect 117 -427 121 -413
rect 145 -427 149 -413
rect 230 -421 234 -413
rect 252 -417 256 -413
rect 95 -443 99 -439
rect 131 -443 135 -431
rect 204 -433 208 -429
rect 216 -437 220 -425
rect 142 -442 158 -438
rect 83 -447 99 -443
rect 106 -447 135 -443
rect -41 -475 -28 -471
rect -15 -475 75 -471
rect -14 -497 -10 -475
rect 8 -497 12 -475
rect 83 -479 87 -447
rect 95 -451 99 -447
rect 109 -471 113 -455
rect 117 -459 121 -447
rect 128 -455 146 -451
rect 145 -471 149 -463
rect 94 -475 95 -471
rect 108 -475 117 -471
rect 121 -475 145 -471
rect 23 -483 87 -479
rect 154 -479 158 -442
rect 194 -441 220 -437
rect 238 -429 242 -421
rect 238 -437 242 -433
rect 277 -429 281 -405
rect 176 -451 180 -441
rect 216 -445 220 -441
rect 165 -455 169 -451
rect 173 -455 180 -451
rect 176 -461 180 -455
rect 187 -457 191 -453
rect 176 -465 193 -461
rect 211 -465 223 -461
rect 230 -471 234 -449
rect 241 -457 245 -453
rect 252 -471 256 -441
rect 185 -475 189 -471
rect 193 -475 202 -471
rect 220 -475 256 -471
rect 277 -479 281 -433
rect 154 -483 277 -479
rect 299 -479 303 -396
rect 313 -405 322 -401
rect 311 -475 322 -471
rect -28 -505 -24 -501
rect -6 -505 -2 -501
rect 23 -502 27 -483
rect 311 -487 318 -475
rect 31 -495 35 -491
rect 41 -491 187 -487
rect 209 -491 216 -487
rect 223 -491 285 -487
rect 295 -491 318 -487
rect -29 -509 -24 -505
rect -17 -509 -2 -505
rect 5 -509 20 -505
rect -28 -513 -24 -509
rect -6 -513 -2 -509
rect 16 -513 31 -509
rect 41 -510 45 -491
rect 209 -495 213 -491
rect 49 -503 53 -499
rect 59 -499 87 -495
rect 94 -499 95 -495
rect 108 -499 154 -495
rect 158 -499 197 -495
rect 208 -499 213 -495
rect 284 -499 288 -491
rect 306 -495 310 -491
rect -14 -535 -10 -517
rect 8 -535 12 -517
rect 16 -517 20 -513
rect 16 -521 49 -517
rect 59 -518 63 -499
rect 67 -511 71 -507
rect 16 -525 20 -521
rect 83 -519 87 -499
rect 109 -511 113 -499
rect 117 -503 121 -499
rect 145 -503 149 -499
rect 201 -503 205 -499
rect 95 -519 99 -515
rect 131 -519 135 -507
rect 142 -518 169 -514
rect 83 -523 99 -519
rect 106 -523 135 -519
rect 187 -519 191 -507
rect 258 -511 262 -507
rect 270 -515 274 -503
rect 248 -519 274 -515
rect 292 -507 296 -499
rect 292 -515 296 -511
rect 198 -523 226 -519
rect 16 -529 67 -525
rect 95 -527 99 -523
rect -41 -539 -28 -535
rect -15 -539 62 -535
rect -41 -542 62 -539
rect 69 -542 79 -535
rect 75 -543 79 -542
rect 109 -543 113 -531
rect 117 -535 121 -523
rect 128 -531 132 -527
rect 145 -543 149 -539
rect 75 -547 95 -543
rect 108 -547 117 -543
rect 121 -547 150 -543
rect 163 -557 167 -531
rect 187 -535 191 -523
rect 222 -529 226 -523
rect 230 -529 234 -519
rect 270 -523 274 -519
rect 222 -533 234 -529
rect 201 -543 205 -539
rect 230 -539 234 -533
rect 241 -535 245 -531
rect 230 -543 247 -539
rect 265 -543 277 -539
rect 175 -547 179 -543
rect 183 -547 187 -543
rect 198 -547 224 -543
rect 220 -549 224 -547
rect 284 -549 288 -527
rect 295 -535 299 -531
rect 306 -535 310 -519
rect 306 -541 322 -535
rect 306 -549 310 -541
rect 220 -553 256 -549
rect 274 -553 322 -549
rect 163 -561 299 -557
rect -41 -569 -21 -562
rect 53 -569 62 -562
rect 69 -566 156 -562
rect 310 -566 322 -562
rect 69 -569 322 -566
rect -17 -584 -13 -569
rect 3 -584 7 -569
rect 23 -584 27 -569
rect 44 -584 48 -569
rect 149 -573 317 -569
rect 55 -580 63 -576
rect -41 -599 -36 -595
rect -41 -607 -36 -603
rect -29 -613 -25 -588
rect -9 -604 -5 -588
rect -18 -608 -5 -604
rect -37 -617 -25 -613
rect -37 -620 -33 -617
rect -29 -620 -25 -617
rect -9 -620 -5 -608
rect 11 -595 15 -588
rect 32 -595 36 -588
rect 52 -595 56 -588
rect 22 -599 36 -595
rect 2 -617 3 -613
rect 11 -620 15 -599
rect 32 -620 36 -599
rect 45 -599 56 -595
rect 62 -595 66 -588
rect 73 -586 77 -580
rect 73 -590 80 -586
rect 62 -599 322 -595
rect 45 -613 49 -599
rect 56 -607 58 -603
rect 62 -607 69 -603
rect 73 -607 322 -603
rect 49 -617 56 -613
rect 52 -620 56 -617
rect 52 -624 63 -620
rect 77 -624 80 -620
rect -17 -630 -13 -624
rect 3 -630 7 -624
rect 23 -630 27 -624
rect 44 -630 48 -624
rect -41 -637 -22 -630
rect 52 -637 216 -630
rect 223 -637 322 -630
rect -41 -638 322 -637
rect -41 -645 60 -638
rect 296 -645 322 -638
rect -33 -654 42 -650
rect 38 -717 42 -654
rect 61 -689 65 -645
rect 88 -681 92 -645
rect 103 -672 107 -666
rect 112 -675 116 -674
rect 112 -681 116 -679
rect 122 -681 126 -645
rect 156 -681 160 -645
rect 77 -700 81 -689
rect 65 -709 68 -705
rect 100 -712 104 -689
rect 146 -703 150 -689
rect 133 -707 146 -703
rect 168 -704 172 -689
rect 175 -691 179 -665
rect 133 -710 137 -707
rect 182 -704 186 -674
rect 199 -691 203 -666
rect 208 -681 212 -645
rect 219 -674 220 -670
rect 235 -681 239 -645
rect 271 -681 275 -678
rect 195 -703 196 -699
rect 208 -709 212 -703
rect 220 -704 224 -689
rect 259 -699 263 -689
rect 278 -695 282 -666
rect 286 -681 290 -645
rect 272 -699 282 -695
rect 298 -692 302 -689
rect 298 -696 313 -692
rect 246 -703 263 -699
rect 224 -708 226 -704
rect 246 -710 250 -703
rect 298 -704 302 -696
rect 271 -709 275 -708
rect 77 -748 81 -716
rect 100 -748 104 -728
rect 122 -748 126 -714
rect 136 -725 140 -721
rect 146 -748 150 -714
rect 168 -748 172 -720
rect 220 -748 224 -720
rect 235 -748 239 -714
rect 249 -725 253 -721
rect 259 -748 263 -714
rect 298 -748 302 -720
rect 309 -736 313 -696
rect -41 -749 322 -748
rect -41 -756 70 -749
rect 306 -756 322 -749
<< metal2 >>
rect -41 218 77 222
rect 81 219 149 222
rect 153 219 173 222
rect 81 218 173 219
rect 177 218 252 222
rect 256 218 322 222
rect 35 179 39 218
rect 90 210 156 214
rect 198 210 249 214
rect 124 177 169 181
rect 204 176 245 180
rect -41 155 110 159
rect 114 155 223 159
rect 227 155 322 159
rect 32 128 43 132
rect 39 53 43 128
rect 39 -72 43 49
rect 61 -20 65 111
rect 112 91 138 95
rect 113 67 155 71
rect 177 -35 181 111
rect 241 53 245 123
rect 262 115 266 144
rect 226 49 256 53
rect 260 49 268 53
rect 71 -56 185 -52
rect 57 -60 75 -56
rect 181 -60 185 -56
rect 105 -69 109 -65
rect 113 -69 117 -65
rect 105 -73 177 -69
rect 173 -75 177 -73
rect 228 -75 232 -73
rect 173 -79 232 -75
rect 30 -92 43 -88
rect 30 -114 34 -92
rect 241 -108 245 49
rect 264 -108 268 49
rect 30 -118 163 -114
rect 159 -126 163 -118
rect -25 -396 223 -392
rect -25 -405 277 -401
rect 281 -405 309 -401
rect 313 -405 322 -401
rect -25 -413 75 -409
rect 75 -471 79 -413
rect -33 -520 -29 -509
rect -33 -524 85 -520
rect 62 -562 69 -542
rect 81 -561 85 -524
rect 117 -543 121 -475
rect 154 -495 158 -413
rect 212 -433 238 -429
rect 281 -433 322 -429
rect 169 -514 173 -455
rect 195 -457 237 -453
rect 189 -479 193 -475
rect 179 -483 193 -479
rect 136 -531 163 -527
rect 179 -543 183 -483
rect 187 -519 191 -491
rect 154 -547 171 -543
rect 80 -566 85 -561
rect 80 -586 84 -566
rect -32 -599 11 -595
rect -32 -607 52 -603
rect 7 -617 45 -613
rect 80 -620 84 -590
rect -37 -650 -33 -624
rect 216 -630 223 -491
rect 266 -511 292 -507
rect 249 -535 291 -531
rect -41 -666 103 -662
rect 107 -665 175 -662
rect 179 -665 199 -662
rect 107 -666 199 -665
rect 203 -666 278 -662
rect 282 -666 322 -662
rect 61 -705 65 -666
rect 116 -674 182 -670
rect 224 -674 275 -670
rect 150 -707 195 -703
rect 230 -708 271 -704
rect -41 -729 136 -725
rect 140 -729 249 -725
rect 253 -729 322 -725
rect 309 -764 313 -740
<< ntransistor >>
rect 51 175 55 177
rect 103 170 105 174
rect 114 170 116 174
rect 177 181 179 185
rect 151 176 153 180
rect 142 171 146 173
rect 194 171 198 173
rect 74 163 78 165
rect 216 170 218 174
rect 227 170 229 174
rect 272 171 276 173
rect 101 83 105 87
rect 123 75 127 79
rect 193 87 197 91
rect 215 87 219 91
rect 163 83 167 87
rect 146 59 150 63
rect 46 -68 50 -64
rect 134 -81 138 -77
rect 84 -95 88 -91
rect 91 -95 95 -91
rect 98 -95 102 -91
rect 120 -95 124 -91
rect 221 -87 225 -83
rect 196 -95 200 -91
rect 203 -95 207 -91
rect 235 -95 239 -91
rect 249 -95 253 -91
rect 54 -100 58 -96
rect 148 -99 152 -95
rect 162 -99 166 -95
rect 31 -506 35 -502
rect 102 -455 106 -451
rect 183 -441 187 -437
rect 124 -463 128 -459
rect 138 -463 142 -459
rect 245 -441 249 -437
rect 223 -449 227 -445
rect 200 -465 204 -461
rect -21 -517 -17 -513
rect 1 -517 5 -513
rect 49 -514 53 -510
rect 67 -522 71 -518
rect 102 -531 106 -527
rect 237 -519 241 -515
rect 124 -539 128 -535
rect 138 -539 142 -535
rect 194 -539 198 -535
rect 299 -519 303 -515
rect 277 -527 281 -523
rect 254 -543 258 -539
rect 69 -580 71 -576
rect -22 -588 -20 -584
rect -2 -588 0 -584
rect 18 -588 20 -584
rect 39 -588 41 -584
rect 58 -588 60 -584
rect 77 -709 81 -707
rect 129 -714 131 -710
rect 140 -714 142 -710
rect 203 -703 205 -699
rect 177 -708 179 -704
rect 168 -713 172 -711
rect 220 -713 224 -711
rect 100 -721 104 -719
rect 242 -714 244 -710
rect 253 -714 255 -710
rect 298 -713 302 -711
<< ptransistor >>
rect 46 195 48 203
rect 69 195 71 203
rect 81 195 83 203
rect 103 195 105 203
rect 114 195 116 203
rect 137 195 139 203
rect 189 195 191 203
rect 216 195 218 203
rect 227 195 229 203
rect 240 195 242 203
rect 267 195 269 203
rect 101 103 105 107
rect 193 103 197 107
rect 215 103 219 107
rect 123 99 127 103
rect 46 -49 50 -45
rect 84 -48 88 -44
rect 91 -48 95 -44
rect 98 -48 102 -44
rect 120 -48 124 -44
rect 148 -48 152 -44
rect 162 -48 166 -44
rect 196 -48 200 -44
rect 203 -48 207 -44
rect 235 -48 239 -44
rect 249 -48 253 -44
rect 54 -84 58 -80
rect 134 -65 138 -61
rect 221 -59 225 -55
rect -21 -501 -17 -497
rect 1 -501 5 -497
rect 245 -421 249 -417
rect 223 -425 227 -421
rect 124 -431 128 -427
rect 138 -431 142 -427
rect 102 -439 106 -435
rect 299 -499 303 -495
rect 277 -503 281 -499
rect 124 -507 128 -503
rect 138 -507 142 -503
rect 194 -507 198 -503
rect 102 -515 106 -511
rect -22 -624 -20 -620
rect -2 -624 0 -620
rect 18 -624 20 -620
rect 39 -624 41 -620
rect 69 -624 71 -620
rect 72 -689 74 -681
rect 95 -689 97 -681
rect 107 -689 109 -681
rect 129 -689 131 -681
rect 140 -689 142 -681
rect 163 -689 165 -681
rect 215 -689 217 -681
rect 242 -689 244 -681
rect 253 -689 255 -681
rect 266 -689 268 -681
rect 293 -689 295 -681
<< polycontact >>
rect -12 239 -4 247
rect 77 208 81 212
rect 189 210 193 214
rect 86 205 90 209
rect 42 175 46 179
rect 124 187 128 191
rect 149 189 153 193
rect 173 189 177 193
rect 182 171 186 175
rect 198 185 202 189
rect 242 185 246 189
rect 110 163 114 167
rect 245 171 249 175
rect 223 163 227 167
rect 123 119 127 123
rect 256 119 260 123
rect 101 91 105 95
rect 193 95 197 99
rect 146 91 150 95
rect 256 100 260 104
rect 215 95 219 99
rect 235 95 239 99
rect 101 67 105 71
rect 163 67 167 71
rect 123 59 127 63
rect -13 49 -5 53
rect 162 41 166 45
rect 84 -23 88 -19
rect 162 -23 166 -19
rect 91 -31 95 -27
rect 148 -31 152 -27
rect 203 -23 207 -19
rect 196 -31 200 -27
rect 235 -31 239 -27
rect 249 -23 253 -19
rect 46 -60 50 -56
rect 54 -92 58 -88
rect 98 -65 102 -61
rect 120 -65 124 -61
rect 134 -73 138 -69
rect 221 -73 225 -69
rect 49 -130 53 -126
rect 31 -139 35 -135
rect 31 -491 35 -487
rect 49 -499 53 -495
rect 67 -147 71 -143
rect -21 -509 -17 -505
rect 1 -509 5 -505
rect 23 -506 27 -502
rect 223 -405 227 -401
rect 245 -405 249 -401
rect 102 -447 106 -443
rect 124 -455 128 -451
rect 200 -433 204 -429
rect 138 -442 142 -438
rect 146 -455 150 -451
rect 161 -455 165 -451
rect 183 -457 187 -453
rect 245 -457 249 -453
rect 223 -465 227 -461
rect 145 -475 149 -471
rect 181 -475 185 -471
rect 277 -483 281 -479
rect 299 -483 303 -479
rect 67 -507 71 -503
rect 41 -514 45 -510
rect 59 -522 63 -518
rect 102 -523 106 -519
rect 124 -531 128 -527
rect 138 -518 142 -514
rect 254 -511 258 -507
rect 194 -523 198 -519
rect 237 -535 241 -531
rect 277 -543 281 -539
rect 299 -535 303 -531
rect 299 -561 303 -557
rect 51 -580 55 -576
rect -22 -608 -18 -604
rect 18 -599 22 -595
rect -2 -617 2 -613
rect 58 -607 62 -603
rect 69 -607 73 -603
rect 103 -676 107 -672
rect 215 -674 219 -670
rect 112 -679 116 -675
rect 68 -709 72 -705
rect 38 -721 42 -717
rect 150 -697 154 -693
rect 175 -695 179 -691
rect 199 -695 203 -691
rect 208 -713 212 -709
rect 224 -699 228 -695
rect 268 -699 272 -695
rect 136 -721 140 -717
rect 271 -713 275 -709
rect 249 -721 253 -717
<< ndcontact >>
rect 51 180 55 184
rect 51 168 55 172
rect 74 168 78 172
rect 96 170 100 174
rect 107 170 111 174
rect 120 170 124 174
rect 170 181 174 185
rect 182 181 186 185
rect 142 176 146 180
rect 156 176 160 180
rect 194 176 198 180
rect 142 164 146 168
rect 209 170 213 174
rect 220 170 224 174
rect 233 170 237 174
rect 272 176 276 180
rect 194 164 198 168
rect 272 164 276 168
rect 74 156 78 160
rect 94 83 98 87
rect 108 83 112 87
rect 116 75 120 79
rect 130 75 134 79
rect 186 87 190 91
rect 200 87 204 91
rect 208 87 212 91
rect 222 87 226 91
rect 156 83 160 87
rect 170 83 174 87
rect 139 59 143 63
rect 153 59 157 63
rect 39 -68 43 -64
rect 53 -68 57 -64
rect 127 -81 131 -77
rect 141 -81 145 -77
rect 77 -95 81 -91
rect 105 -95 109 -91
rect 113 -95 117 -91
rect 127 -95 131 -91
rect 214 -87 218 -83
rect 228 -87 232 -83
rect 189 -95 193 -91
rect 210 -95 214 -91
rect 228 -95 232 -91
rect 242 -95 246 -91
rect 256 -95 260 -91
rect 47 -100 51 -96
rect 61 -100 65 -96
rect 140 -99 144 -95
rect 155 -99 159 -95
rect 169 -99 173 -95
rect 31 -499 35 -495
rect 95 -455 99 -451
rect 109 -455 113 -451
rect 176 -441 180 -437
rect 190 -441 194 -437
rect 117 -463 121 -459
rect 145 -463 149 -459
rect 238 -441 242 -437
rect 252 -441 256 -437
rect 216 -449 220 -445
rect 230 -449 234 -445
rect 193 -465 197 -461
rect 207 -465 211 -461
rect 31 -513 35 -509
rect 49 -507 53 -503
rect -28 -517 -24 -513
rect -14 -517 -10 -513
rect -6 -517 -2 -513
rect 8 -517 12 -513
rect 49 -521 53 -517
rect 67 -515 71 -511
rect 67 -529 71 -525
rect 95 -531 99 -527
rect 109 -531 113 -527
rect 230 -519 234 -515
rect 244 -519 248 -515
rect 117 -539 121 -535
rect 145 -539 149 -535
rect 187 -539 191 -535
rect 201 -539 205 -535
rect 292 -519 296 -515
rect 306 -519 310 -515
rect 270 -527 274 -523
rect 284 -527 288 -523
rect 247 -543 251 -539
rect 261 -543 265 -539
rect 63 -580 67 -576
rect 73 -580 77 -576
rect -29 -588 -25 -584
rect -17 -588 -13 -584
rect -9 -588 -5 -584
rect 3 -588 7 -584
rect 11 -588 15 -584
rect 23 -588 27 -584
rect 32 -588 36 -584
rect 44 -588 48 -584
rect 52 -588 56 -584
rect 62 -588 66 -584
rect 77 -704 81 -700
rect 77 -716 81 -712
rect 100 -716 104 -712
rect 122 -714 126 -710
rect 133 -714 137 -710
rect 146 -714 150 -710
rect 196 -703 200 -699
rect 208 -703 212 -699
rect 168 -708 172 -704
rect 182 -708 186 -704
rect 220 -708 224 -704
rect 168 -720 172 -716
rect 235 -714 239 -710
rect 246 -714 250 -710
rect 259 -714 263 -710
rect 298 -708 302 -704
rect 220 -720 224 -716
rect 298 -720 302 -716
rect 100 -728 104 -724
<< pdcontact >>
rect 39 195 43 203
rect 51 195 55 203
rect 62 195 66 203
rect 74 195 78 203
rect 86 195 90 203
rect 96 195 100 203
rect 120 195 124 203
rect 130 195 134 203
rect 142 195 146 203
rect 182 195 186 203
rect 194 195 198 203
rect 209 195 213 203
rect 233 195 237 203
rect 245 195 249 203
rect 260 195 264 203
rect 272 195 276 203
rect 94 103 98 107
rect 108 103 112 107
rect 186 103 190 107
rect 200 103 204 107
rect 208 103 212 107
rect 222 103 226 107
rect 116 99 120 103
rect 130 99 134 103
rect 39 -49 43 -45
rect 53 -49 57 -45
rect 77 -48 81 -44
rect 105 -48 109 -44
rect 113 -48 117 -44
rect 128 -48 132 -44
rect 140 -48 144 -44
rect 155 -48 159 -44
rect 169 -48 173 -44
rect 189 -48 193 -44
rect 210 -48 214 -44
rect 228 -48 232 -44
rect 242 -48 246 -44
rect 256 -48 260 -44
rect 47 -84 51 -80
rect 61 -84 65 -80
rect 127 -65 131 -61
rect 141 -65 145 -61
rect 214 -59 218 -55
rect 228 -59 232 -55
rect -28 -501 -24 -497
rect -14 -501 -10 -497
rect -6 -501 -2 -497
rect 8 -501 12 -497
rect 238 -421 242 -417
rect 252 -421 256 -417
rect 216 -425 220 -421
rect 230 -425 234 -421
rect 117 -431 121 -427
rect 131 -431 135 -427
rect 145 -431 149 -427
rect 95 -439 99 -435
rect 109 -439 113 -435
rect 292 -499 296 -495
rect 306 -499 310 -495
rect 270 -503 274 -499
rect 284 -503 288 -499
rect 117 -507 121 -503
rect 131 -507 135 -503
rect 145 -507 149 -503
rect 187 -507 191 -503
rect 201 -507 205 -503
rect 95 -515 99 -511
rect 109 -515 113 -511
rect -29 -624 -25 -620
rect -17 -624 -13 -620
rect -9 -624 -5 -620
rect 3 -624 7 -620
rect 11 -624 15 -620
rect 23 -624 27 -620
rect 32 -624 36 -620
rect 44 -624 48 -620
rect 63 -624 67 -620
rect 73 -624 77 -620
rect 65 -689 69 -681
rect 77 -689 81 -681
rect 88 -689 92 -681
rect 100 -689 104 -681
rect 112 -689 116 -681
rect 122 -689 126 -681
rect 146 -689 150 -681
rect 156 -689 160 -681
rect 168 -689 172 -681
rect 208 -689 212 -681
rect 220 -689 224 -681
rect 235 -689 239 -681
rect 259 -689 263 -681
rect 271 -689 275 -681
rect 286 -689 290 -681
rect 298 -689 302 -681
<< m2contact >>
rect 77 218 81 222
rect 86 210 90 214
rect 149 219 153 223
rect 35 175 39 179
rect 120 177 124 181
rect 173 218 177 222
rect 156 210 160 214
rect 194 210 198 214
rect 252 218 256 222
rect 245 206 249 210
rect 165 181 169 185
rect 200 176 204 180
rect 245 176 249 180
rect 110 155 114 159
rect 223 155 227 159
rect 262 144 266 148
rect 19 128 32 136
rect 61 111 65 115
rect 177 111 181 115
rect 262 111 266 115
rect 108 91 112 95
rect 138 91 142 95
rect 109 67 113 71
rect 155 67 159 71
rect 256 74 260 78
rect 39 49 43 53
rect 222 49 226 53
rect 61 -24 65 -20
rect 177 -39 181 -35
rect 53 -60 57 -56
rect 39 -76 43 -72
rect 105 -65 109 -61
rect 113 -65 117 -61
rect 181 -64 185 -60
rect 228 -73 232 -69
rect 256 -73 260 -69
rect 43 -92 47 -88
rect 241 -112 245 -108
rect 264 -112 268 -108
rect 159 -130 163 -126
rect -29 -396 -25 -392
rect 223 -396 227 -392
rect -29 -405 -25 -401
rect 277 -405 281 -401
rect -29 -413 -25 -409
rect 75 -413 79 -409
rect 154 -413 158 -409
rect 208 -433 212 -429
rect 75 -475 79 -471
rect 117 -475 121 -471
rect 238 -433 242 -429
rect 277 -433 281 -429
rect 169 -455 173 -451
rect 191 -457 195 -453
rect 237 -457 241 -453
rect 189 -475 193 -471
rect 309 -405 313 -401
rect 187 -491 191 -487
rect 216 -491 223 -487
rect -33 -509 -29 -505
rect 154 -499 158 -495
rect 169 -518 173 -514
rect 262 -511 266 -507
rect 292 -511 296 -507
rect 187 -523 191 -519
rect 62 -542 69 -535
rect 132 -531 136 -527
rect 163 -531 167 -527
rect 117 -547 121 -543
rect 150 -547 154 -543
rect 245 -535 249 -531
rect 171 -547 175 -543
rect 179 -547 183 -543
rect 291 -535 295 -531
rect 62 -569 69 -562
rect -36 -599 -32 -595
rect -36 -607 -32 -603
rect -37 -624 -33 -620
rect 11 -599 15 -595
rect 3 -617 7 -613
rect 80 -590 84 -586
rect 52 -607 56 -603
rect 45 -617 49 -613
rect 80 -624 84 -620
rect 216 -637 223 -630
rect -37 -654 -33 -650
rect 103 -666 107 -662
rect 112 -674 116 -670
rect 175 -665 179 -661
rect 61 -709 65 -705
rect 146 -707 150 -703
rect 199 -666 203 -662
rect 182 -674 186 -670
rect 220 -674 224 -670
rect 278 -666 282 -662
rect 271 -678 275 -674
rect 191 -703 195 -699
rect 226 -708 230 -704
rect 271 -708 275 -704
rect 136 -729 140 -725
rect 249 -729 253 -725
rect 309 -740 313 -736
<< psubstratepcontact >>
rect 44 128 280 135
rect 98 49 116 53
rect 61 -69 65 -63
rect 117 -112 134 -108
rect 95 -475 108 -471
rect 202 -475 220 -471
rect -28 -539 -15 -535
rect 95 -547 108 -543
rect 187 -547 198 -543
rect 256 -553 274 -549
rect -21 -569 53 -562
rect 70 -756 306 -749
<< nsubstratencontact >>
rect 34 239 270 246
rect 109 111 119 115
rect 117 -39 134 -35
rect 36 -85 40 -79
rect -28 -475 -15 -471
rect 95 -413 108 -409
rect 231 -413 241 -409
rect 95 -499 108 -495
rect 197 -499 208 -495
rect 285 -491 295 -487
rect -22 -637 52 -630
rect 60 -645 296 -638
<< labels >>
rlabel metal1 37 92 37 92 1 kris_bit_1_0/Qout
rlabel metal2 -32 -521 -31 -521 3 kris_bit_1_0/shiftbit_in
rlabel metal2 309 -764 313 -764 1 kris_bit_1_0/regout
rlabel metal1 272 184 276 188 3 kris_bit_1_0/reg2_na_0/Qout
rlabel metal1 54 239 57 247 7 kris_bit_1_0/reg2_na_0/Vdd
rlabel metal1 55 128 59 136 7 kris_bit_1_0/reg2_na_0/GND
rlabel metal2 33 218 37 222 7 kris_bit_1_0/reg2_na_0/clk
rlabel metal2 39 155 43 159 7 kris_bit_1_0/reg2_na_0/rst
rlabel polysilicon 38 163 42 165 7 kris_bit_1_0/reg2_na_0/Din
rlabel polysilicon 103 122 103 122 5 kris_bit_1_0/add1_flat_first_0/B
rlabel metal1 72 114 72 114 5 kris_bit_1_0/add1_flat_first_0/Vdd
rlabel metal1 133 50 133 50 1 kris_bit_1_0/add1_flat_first_0/GND
rlabel metal1 133 114 133 114 5 kris_bit_1_0/add1_flat_first_0/Vdd
rlabel metal1 177 71 177 71 7 kris_bit_1_0/add1_flat_first_0/Out
rlabel metal1 30 -39 30 -35 7 kris_bit_1_0/add1_flat_first_0/Vdd
rlabel polysilicon 237 -17 237 -17 1 kris_bit_1_0/add1_flat_first_0/B
rlabel polysilicon 164 -16 164 -16 5 kris_bit_1_0/add1_flat_first_0/A
rlabel metal1 163 -36 163 -36 5 kris_bit_1_0/add1_flat_first_0/Vdd
rlabel metal1 163 -111 163 -111 1 kris_bit_1_0/add1_flat_first_0/GND
rlabel metal1 36 -58 36 -58 3 kris_bit_1_0/add1_flat_first_0/Cout
rlabel metal1 32 -58 32 -58 3 kris_bit_1_0/add1_flat_first_0/Cout
rlabel metal1 261 -111 261 -111 1 kris_bit_1_0/add1_flat_first_0/GND
rlabel metal1 133 43 133 43 1 kris_bit_1_0/add1_flat_first_0/a0
rlabel metal1 133 35 133 35 1 kris_bit_1_0/add1_flat_first_0/a1
rlabel metal1 133 27 133 27 1 kris_bit_1_0/add1_flat_first_0/a2
rlabel metal1 133 19 133 19 1 kris_bit_1_0/add1_flat_first_0/a3
rlabel metal1 133 11 133 11 1 kris_bit_1_0/add1_flat_first_0/a4
rlabel metal1 133 2 133 2 1 kris_bit_1_0/add1_flat_first_0/a5
rlabel metal1 133 -5 133 -5 1 kris_bit_1_0/add1_flat_first_0/a6
rlabel metal1 133 -13 133 -13 1 kris_bit_1_0/add1_flat_first_0/a6
rlabel metal1 267 -71 267 -71 7 kris_bit_1_0/add1_flat_first_0/Cin
rlabel metal1 263 -71 263 -71 7 kris_bit_1_0/add1_flat_first_0/Cin
rlabel metal2 161 -125 161 -125 1 kris_bit_1_0/add1_flat_first_0/S
rlabel metal2 161 -121 161 -121 1 kris_bit_1_0/add1_flat_first_0/S
rlabel metal1 86 -410 86 -410 5 kris_bit_1_0/mux1_0/Vdd
rlabel metal1 82 -546 82 -546 1 kris_bit_1_0/mux1_0/GND
rlabel polysilicon 33 -464 33 -464 5 kris_bit_1_0/mux1_0/In0
rlabel polysilicon 51 -464 51 -464 5 kris_bit_1_0/mux1_0/In1
rlabel polysilicon 69 -464 69 -464 5 kris_bit_1_0/mux1_0/In2
rlabel metal1 -39 -411 -39 -411 3 kris_bit_1_0/mux1_0/Vdd
rlabel metal1 -39 -403 -39 -403 3 kris_bit_1_0/mux1_0/sel0
rlabel metal1 -39 -394 -39 -394 3 kris_bit_1_0/mux1_0/sel1
rlabel metal1 105 -201 105 -201 1 kris_bit_1_0/mux1_0/zero
rlabel metal1 99 -264 99 -264 1 kris_bit_1_0/mux1_0/rbit0
rlabel metal1 99 -257 99 -257 1 kris_bit_1_0/mux1_0/zero
rlabel metal1 99 -248 99 -248 1 kris_bit_1_0/mux1_0/zero
rlabel metal1 99 -240 99 -240 1 kris_bit_1_0/mux1_0/zero
rlabel metal1 99 -233 99 -233 1 kris_bit_1_0/mux1_0/zero
rlabel metal1 99 -224 99 -224 1 kris_bit_1_0/mux1_0/zero
rlabel metal1 99 -216 99 -216 1 kris_bit_1_0/mux1_0/zero
rlabel metal1 98 -208 98 -208 1 kris_bit_1_0/mux1_0/zero
rlabel metal1 97 -191 97 -191 1 kris_bit_1_0/mux1_0/dvdin7
rlabel metal1 97 -184 97 -184 1 kris_bit_1_0/mux1_0/dvdin6
rlabel metal1 96 -176 96 -176 1 kris_bit_1_0/mux1_0/dvdin5
rlabel metal1 96 -168 96 -168 1 kris_bit_1_0/mux1_0/dvdin4
rlabel metal1 96 -160 96 -160 1 kris_bit_1_0/mux1_0/dvdin3
rlabel metal1 96 -153 96 -153 1 kris_bit_1_0/mux1_0/dvdin2
rlabel metal1 96 -145 96 -145 1 kris_bit_1_0/mux1_0/dvdin1
rlabel metal1 96 -137 96 -137 1 kris_bit_1_0/mux1_0/dvdin0
rlabel metal1 99 -272 99 -272 1 kris_bit_1_0/mux1_0/rbi1
rlabel metal1 99 -281 99 -281 1 kris_bit_1_0/mux1_0/rbit2
rlabel metal1 98 -288 98 -288 1 kris_bit_1_0/mux1_0/rbit3
rlabel metal1 99 -295 99 -295 1 kris_bit_1_0/mux1_0/rbit4
rlabel metal1 99 -303 99 -303 1 kris_bit_1_0/mux1_0/rbit5
rlabel metal1 98 -310 98 -310 1 kris_bit_1_0/mux1_0/rbit6
rlabel metal1 99 -319 99 -319 1 kris_bit_1_0/mux1_0/rbit7
rlabel metal1 98 -327 98 -327 1 kris_bit_1_0/mux1_0/rbit8
rlabel metal1 99 -335 99 -335 1 kris_bit_1_0/mux1_0/rbit9
rlabel metal1 98 -343 98 -343 1 kris_bit_1_0/mux1_0/rbit10
rlabel metal1 98 -351 98 -351 1 kris_bit_1_0/mux1_0/rbit11
rlabel metal1 99 -359 99 -359 1 kris_bit_1_0/mux1_0/rbit12
rlabel metal1 99 -367 99 -367 1 kris_bit_1_0/mux1_0/rbit13
rlabel metal1 98 -375 98 -375 1 kris_bit_1_0/mux1_0/rbit14
rlabel metal1 98 -384 98 -384 1 kris_bit_1_0/mux1_0/rbit15
rlabel metal1 78 -481 78 -481 7 kris_bit_1_0/mux1_0/31MUX_0/Sel0
rlabel metal1 78 -489 78 -489 7 kris_bit_1_0/mux1_0/31MUX_0/Sel1
rlabel metal1 78 -497 78 -497 7 kris_bit_1_0/mux1_0/31MUX_0/Sel2
rlabel polysilicon 33 -468 33 -468 5 kris_bit_1_0/mux1_0/31MUX_0/In0
rlabel polysilicon 51 -468 51 -468 5 kris_bit_1_0/mux1_0/31MUX_0/In1
rlabel polysilicon 69 -468 69 -468 5 kris_bit_1_0/mux1_0/31MUX_0/In2
rlabel metal1 10 -538 10 -538 1 kris_bit_1_0/mux1_0/31MUX_0/GND
rlabel metal1 -31 -507 -31 -507 3 kris_bit_1_0/mux1_0/31MUX_0/Out
rlabel metal1 10 -472 10 -472 5 kris_bit_1_0/mux1_0/31MUX_0/Vdd
rlabel metal1 88 -489 88 -489 3 kris_bit_1_0/mux1_0/MUXsel_0/Out00
rlabel metal1 162 -410 162 -410 5 kris_bit_1_0/mux1_0/MUXsel_0/Vdd
rlabel metal1 161 -496 161 -496 5 kris_bit_1_0/mux1_0/MUXsel_0/Vdd
rlabel metal1 88 -445 88 -445 3 kris_bit_1_0/mux1_0/MUXsel_0/Out10
rlabel metal1 88 -521 88 -521 3 kris_bit_1_0/mux1_0/MUXsel_0/Out01
rlabel metal1 179 -546 179 -546 1 kris_bit_1_0/mux1_0/MUXsel_0/GND
rlabel metal2 321 -431 321 -431 7 kris_bit_1_0/mux1_0/MUXsel_0/Sel0
rlabel metal1 322 -405 322 -401 7 kris_bit_1_0/mux1_0/MUXsel_0/sel0
rlabel metal1 322 -396 322 -392 6 kris_bit_1_0/mux1_0/MUXsel_0/sel1
rlabel psubstratepcontact 217 -474 217 -474 1 kris_bit_1_0/mux1_0/MUXsel_0/XOR_0/GND
rlabel metal1 217 -410 217 -410 5 kris_bit_1_0/mux1_0/MUXsel_0/XOR_0/Vdd
rlabel polysilicon 247 -406 247 -406 5 kris_bit_1_0/mux1_0/MUXsel_0/XOR_0/In1
rlabel polysilicon 225 -406 225 -406 5 kris_bit_1_0/mux1_0/MUXsel_0/XOR_0/In2
rlabel metal1 173 -453 173 -453 3 kris_bit_1_0/mux1_0/MUXsel_0/XOR_0/Out
rlabel psubstratepcontact 271 -552 271 -552 1 kris_bit_1_0/mux1_0/MUXsel_0/XOR_1/GND
rlabel metal1 271 -488 271 -488 5 kris_bit_1_0/mux1_0/MUXsel_0/XOR_1/Vdd
rlabel polysilicon 301 -484 301 -484 5 kris_bit_1_0/mux1_0/MUXsel_0/XOR_1/In1
rlabel polysilicon 279 -484 279 -484 5 kris_bit_1_0/mux1_0/MUXsel_0/XOR_1/In2
rlabel metal1 227 -531 227 -531 3 kris_bit_1_0/mux1_0/MUXsel_0/XOR_1/Out
rlabel metal1 78 -599 90 -595 3 kris_bit_1_0/shift1_0/inbit
rlabel metal1 78 -607 90 -603 3 kris_bit_1_0/shift1_0/shift
rlabel metal1 -41 -599 -34 -595 7 kris_bit_1_0/shift1_0/inbit_next
rlabel metal1 -41 -607 -32 -603 7 kris_bit_1_0/shift1_0/shift
rlabel metal2 80 -561 84 -561 1 kris_bit_1_0/shift1_0/shiftbit_in
rlabel metal2 -37 -638 -33 -638 5 kris_bit_1_0/shift1_0/shiftbit_out
rlabel metal1 81 -633 81 -633 1 kris_bit_1_0/shift1_0/Vdd
rlabel metal1 78 -565 78 -565 5 kris_bit_1_0/shift1_0/GND
rlabel metal1 298 -700 302 -696 3 kris_bit_1_0/reg2_na_1/Qout
rlabel metal1 80 -645 83 -637 7 kris_bit_1_0/reg2_na_1/Vdd
rlabel metal1 81 -756 85 -748 7 kris_bit_1_0/reg2_na_1/GND
rlabel metal2 59 -666 63 -662 7 kris_bit_1_0/reg2_na_1/clk
rlabel metal2 65 -729 69 -725 7 kris_bit_1_0/reg2_na_1/rst
rlabel polysilicon 64 -721 68 -719 7 kris_bit_1_0/reg2_na_1/Din
<< end >>
