magic
tech scmos
timestamp 1385599424
<< error_s >>
rect 219 150 224 154
<< polysilicon >>
rect -56 88 -52 420
rect -38 80 -34 429
rect -20 79 -16 420
<< metal1 >>
rect -118 674 40 678
rect -118 666 38 670
rect -127 416 275 420
rect -127 408 275 412
rect -127 400 275 404
rect -127 393 275 397
rect -127 385 275 389
rect -127 377 275 381
rect -127 369 275 373
rect -127 361 275 365
rect -127 353 275 357
rect -127 345 275 349
rect -127 337 275 341
rect -127 329 275 333
rect -127 321 275 325
rect -127 313 275 317
rect -127 305 275 309
rect -127 297 275 301
rect -127 289 275 293
rect -127 281 275 285
rect -127 273 275 277
rect -127 266 275 270
rect -127 258 275 262
rect -127 250 275 254
rect -127 242 275 246
rect -127 234 275 238
rect -127 226 275 230
rect -127 218 275 222
rect -127 210 275 214
rect -127 202 275 206
rect -127 194 275 198
rect -127 186 275 190
rect -127 178 275 182
rect -127 170 275 174
rect -127 159 -116 163
rect -127 150 -116 154
rect -127 142 -116 146
rect -8 142 7 146
rect -4 76 0 112
rect -14 72 0 76
rect -14 64 0 68
rect -14 56 0 60
rect -127 46 -115 50
rect -4 32 0 56
rect -12 12 -8 20
rect -12 8 7 12
<< metal2 >>
rect -112 159 136 163
rect -112 150 222 154
rect 226 150 235 154
rect -112 142 -12 146
rect -12 84 -8 142
<< m2contact >>
rect -116 159 -112 163
rect 136 159 140 163
rect -116 150 -112 154
rect 222 150 226 154
rect -116 142 -112 146
rect -12 142 -8 146
rect -12 80 -8 84
use 31MUX  31MUX_0
timestamp 1385597075
transform 1 0 -61 0 1 58
box -58 -43 53 30
use MUXsel  MUXsel_0
timestamp 1385597418
transform 1 0 157 0 1 204
box -157 -210 78 -41
<< labels >>
rlabel metal1 -1 145 -1 145 5 Vdd
rlabel metal1 -5 9 -5 9 1 GND
rlabel polysilicon -54 91 -54 91 5 In0
rlabel polysilicon -36 91 -36 91 5 In1
rlabel polysilicon -18 91 -18 91 5 In2
rlabel metal1 -126 144 -126 144 3 Vdd
rlabel metal1 -126 152 -126 152 3 sel0
rlabel metal1 -126 161 -126 161 3 sel1
rlabel metal1 -127 416 275 420 5 dvdin0
rlabel metal1 -127 408 275 412 1 dvdin1
rlabel metal1 -127 400 275 404 1 dvdin2
rlabel metal1 -127 393 275 397 1 dvdin3
rlabel metal1 -127 385 275 389 1 dvdin4
rlabel metal1 -127 377 275 381 1 dvdin5
rlabel metal1 -127 369 275 373 1 dvdin6
rlabel metal1 -127 361 275 365 1 dvdin7
rlabel metal1 -127 345 275 349 1 zero
rlabel metal1 -127 353 275 357 1 zero
rlabel metal1 -127 337 275 341 1 zero
rlabel metal1 -127 329 275 333 1 zero
rlabel metal1 -127 321 275 325 1 zero
rlabel metal1 -127 313 275 317 1 zero
rlabel metal1 -127 305 275 309 1 zero
rlabel metal1 -127 297 275 301 1 zero
rlabel metal1 -127 281 275 285 1 rbit1
rlabel metal1 -127 289 275 293 1 rbit0
rlabel metal1 -127 273 275 277 1 rbit2
rlabel metal1 -127 266 275 270 1 rbit3
rlabel metal1 -127 258 275 262 1 rbit4
rlabel metal1 -127 250 275 254 1 rbit5
rlabel metal1 -127 234 275 238 1 rbit7
rlabel metal1 -127 242 275 246 1 rbit6
rlabel metal1 -127 226 275 230 1 rbit8
rlabel metal1 -127 218 275 222 1 rbit9
rlabel metal1 -127 210 275 214 1 rbit10
rlabel metal1 -127 202 275 206 1 rbit11
rlabel metal1 -127 194 275 198 1 rbit12
rlabel metal1 -127 186 275 190 1 rbit13
rlabel metal1 -127 178 275 182 1 rbit14
rlabel metal1 -127 170 275 174 1 rbit15
<< end >>
