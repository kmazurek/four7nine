magic
tech scmos
timestamp 1385162186
<< pwell >>
rect -67 -23 -47 -7
rect -67 -39 75 -23
<< nwell >>
rect -67 -3 75 19
rect -43 -13 75 -3
<< polysilicon >>
rect -59 8 -55 22
rect -59 -8 -55 4
rect -31 -8 -27 22
rect -3 8 1 10
rect 11 8 15 22
rect 33 8 37 10
rect -3 0 1 4
rect -59 -14 -55 -12
rect -31 -24 -27 -12
rect -3 -24 1 -4
rect 11 -24 15 4
rect 33 -16 37 4
rect 63 -8 67 -6
rect 33 -24 37 -20
rect 63 -16 67 -12
rect 63 -24 67 -20
rect -31 -30 -27 -28
rect -3 -30 1 -28
rect 11 -30 15 -28
rect 33 -30 37 -28
rect 63 -30 67 -28
<< ndiffusion >>
rect -62 -12 -59 -8
rect -55 -12 -52 -8
rect -34 -28 -31 -24
rect -27 -28 -24 -24
rect -6 -28 -3 -24
rect 1 -28 11 -24
rect 15 -28 33 -24
rect 37 -28 40 -24
rect 60 -28 63 -24
rect 67 -28 70 -24
<< pdiffusion >>
rect -62 4 -59 8
rect -55 4 -52 8
rect -6 4 -3 8
rect 1 4 4 8
rect 8 4 11 8
rect 15 4 18 8
rect 30 4 33 8
rect 37 4 40 8
rect -34 -12 -31 -8
rect -27 -12 -24 -8
rect 60 -12 63 -8
rect 67 -12 70 -8
<< metal1 >>
rect -66 14 -51 18
rect -38 14 74 18
rect -66 8 -62 14
rect -52 0 -48 4
rect -52 -8 -48 -4
rect -38 -8 -34 14
rect -10 8 -6 14
rect 18 8 22 14
rect 40 8 44 14
rect -6 -4 -3 0
rect 4 -6 8 4
rect 26 -6 30 4
rect 4 -10 52 -6
rect -66 -34 -62 -12
rect -24 -16 -20 -12
rect -24 -20 33 -16
rect -24 -24 -20 -20
rect 40 -24 44 -10
rect 48 -16 52 -10
rect 56 -8 60 14
rect 70 -16 74 -12
rect 48 -20 63 -16
rect 70 -20 78 -16
rect 70 -24 74 -20
rect -38 -34 -34 -28
rect -10 -34 -6 -28
rect 56 -34 60 -28
rect -66 -38 -51 -34
rect -38 -38 74 -34
<< metal2 >>
rect -48 -4 -10 0
<< ntransistor >>
rect -59 -12 -55 -8
rect -31 -28 -27 -24
rect -3 -28 1 -24
rect 11 -28 15 -24
rect 33 -28 37 -24
rect 63 -28 67 -24
<< ptransistor >>
rect -59 4 -55 8
rect -3 4 1 8
rect 11 4 15 8
rect 33 4 37 8
rect -31 -12 -27 -8
rect 63 -12 67 -8
<< polycontact >>
rect -3 -4 1 0
rect 33 -20 37 -16
rect 63 -20 67 -16
<< ndcontact >>
rect -66 -12 -62 -8
rect -52 -12 -48 -8
rect -38 -28 -34 -24
rect -24 -28 -20 -24
rect -10 -28 -6 -24
rect 40 -28 44 -24
rect 56 -28 60 -24
rect 70 -28 74 -24
<< pdcontact >>
rect -66 4 -62 8
rect -52 4 -48 8
rect -10 4 -6 8
rect 4 4 8 8
rect 18 4 22 8
rect 26 4 30 8
rect 40 4 44 8
rect -38 -12 -34 -8
rect -24 -12 -20 -8
rect 56 -12 60 -8
rect 70 -12 74 -8
<< m2contact >>
rect -52 -4 -48 0
rect -10 -4 -6 0
<< psubstratepcontact >>
rect -51 -38 -38 -34
<< nsubstratencontact >>
rect -51 14 -38 18
<< labels >>
rlabel metal1 -8 17 -8 17 5 Vdd
rlabel metal1 -8 -37 -8 -37 1 GND
rlabel polysilicon -57 21 -57 21 5 y1
rlabel polysilicon -29 21 -29 21 5 t
rlabel polysilicon 13 21 13 21 5 y0
rlabel metal1 77 -18 77 -18 7 OutY1
<< end >>
